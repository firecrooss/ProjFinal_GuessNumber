----------------------------------------------------------------------------------------------------------------------------------------------------------------
-- LSD.TOS, April 2018 (DO NOT REMOVE THIS LINE), VHDL 2008
--
-- Pseudo-random number generator.
--
-- This entity has two architectures:
--   heavy ... perhaps better at generating pseudo-random numbers, but uses more configurable logic elements and gives rise to a longer compilation time
--   basic ... weaker pseudo-random number generator (but perfectly acceptable for most purposes)
-- Warning: do not use the rnd output in the very first 10 or so clock cycles (may not be random enough).
--
-- While developing a project that uses this entity keep in mind the following:
-- * two or more instantiations of the pseudo-random number generator require either different architectures of different seed values,
-- * it is better to leave a generator always running (enable always at '1') and to use the pseudo-random number at the times when it is needed; in
--   particular, if the time when the pseudo-random number is used is the result of a key of the kit being pressed, then the number would be truly random
--
-- A simple example of the use of the pseudo_random_generator entity can be found in the file pseudo_random_generator_example_tl.vhd
--

library IEEE;
use     IEEE.STD_LOGIC_1164.ALL;
use     IEEE.NUMERIC_STD.ALL;

entity pseudo_random_generator is
  generic
  (
    N_BITS : integer range 1 to 24 := 18;        -- number of pseudo-random output bits
    SEED   : std_logic_vector(47 downto 0) := "011011101001011011011010011011101001011011011010" -- initial state of the generator
  );
  port
  (
    clock  : in  std_logic;                          -- main clock
    enable : in  std_logic := '1';                   -- when active, the generator produces a new pseudo-random number
    rnd    : out std_logic_vector(N_BITS-1 downto 0) -- pseudo-random bits
  );
end pseudo_random_generator;

--
-- Multi-stage substitution-permutation network (period=2^48, data generated by c_code/pseudo_random_generator.c with n=48 and seed=1)
--
architecture heavy of pseudo_random_generator is
  signal carry    : std_logic := '0';                      -- carry signal between the two halves of the counter
  signal state_00 : std_logic_vector(47 downto 0) := SEED; -- the pseudo-random generator internal counter
  -- state 1 and all relevant data to update it
  signal state_01 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #1
  signal addr_00x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_01_00 : std_logic_vector(15 downto 0) := "0011010101011010";
  constant S_BOX_01_01 : std_logic_vector(15 downto 0) := "0000111100111001";
  constant S_BOX_01_02 : std_logic_vector(15 downto 0) := "0110001100010111";
  constant S_BOX_01_03 : std_logic_vector(15 downto 0) := "1010011101100100";
  signal addr_00x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_01_04 : std_logic_vector(15 downto 0) := "1000101011001110";
  constant S_BOX_01_05 : std_logic_vector(15 downto 0) := "0001110111000101";
  constant S_BOX_01_06 : std_logic_vector(15 downto 0) := "1011011001010100";
  constant S_BOX_01_07 : std_logic_vector(15 downto 0) := "0001001011110011";
  signal addr_00x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_01_08 : std_logic_vector(15 downto 0) := "1001101010011001";
  constant S_BOX_01_09 : std_logic_vector(15 downto 0) := "0000101001110111";
  constant S_BOX_01_10 : std_logic_vector(15 downto 0) := "0000011111011010";
  constant S_BOX_01_11 : std_logic_vector(15 downto 0) := "1010101100001110";
  signal addr_00x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_01_12 : std_logic_vector(15 downto 0) := "1100011100101100";
  constant S_BOX_01_13 : std_logic_vector(15 downto 0) := "1111010100010010";
  constant S_BOX_01_14 : std_logic_vector(15 downto 0) := "0100111001110010";
  constant S_BOX_01_15 : std_logic_vector(15 downto 0) := "0010010111111000";
  signal addr_00x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_01_16 : std_logic_vector(15 downto 0) := "1001010010101101";
  constant S_BOX_01_17 : std_logic_vector(15 downto 0) := "1100110001011100";
  constant S_BOX_01_18 : std_logic_vector(15 downto 0) := "1001110111000010";
  constant S_BOX_01_19 : std_logic_vector(15 downto 0) := "1011000001010111";
  signal addr_00x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_01_20 : std_logic_vector(15 downto 0) := "0001011000111011";
  constant S_BOX_01_21 : std_logic_vector(15 downto 0) := "1010011011100010";
  constant S_BOX_01_22 : std_logic_vector(15 downto 0) := "1111000000100111";
  constant S_BOX_01_23 : std_logic_vector(15 downto 0) := "0010110010001111";
  signal addr_00x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_01_24 : std_logic_vector(15 downto 0) := "1100111010001001";
  constant S_BOX_01_25 : std_logic_vector(15 downto 0) := "0111000011101001";
  constant S_BOX_01_26 : std_logic_vector(15 downto 0) := "0010110101001011";
  constant S_BOX_01_27 : std_logic_vector(15 downto 0) := "1111100100010001";
  signal addr_00x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_01_28 : std_logic_vector(15 downto 0) := "0101001011001011";
  constant S_BOX_01_29 : std_logic_vector(15 downto 0) := "0100011100010111";
  constant S_BOX_01_30 : std_logic_vector(15 downto 0) := "1000110011010011";
  constant S_BOX_01_31 : std_logic_vector(15 downto 0) := "0110110110001001";
  signal addr_00x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_01_32 : std_logic_vector(15 downto 0) := "1111100010000011";
  constant S_BOX_01_33 : std_logic_vector(15 downto 0) := "0110001100101011";
  constant S_BOX_01_34 : std_logic_vector(15 downto 0) := "1000100101011011";
  constant S_BOX_01_35 : std_logic_vector(15 downto 0) := "1101010000111001";
  signal addr_00x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_01_36 : std_logic_vector(15 downto 0) := "0011000110001111";
  constant S_BOX_01_37 : std_logic_vector(15 downto 0) := "0011110011100010";
  constant S_BOX_01_38 : std_logic_vector(15 downto 0) := "1110010100101010";
  constant S_BOX_01_39 : std_logic_vector(15 downto 0) := "1010001011101001";
  signal addr_00x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_01_40 : std_logic_vector(15 downto 0) := "1000111000101101";
  constant S_BOX_01_41 : std_logic_vector(15 downto 0) := "0010101111101000";
  constant S_BOX_01_42 : std_logic_vector(15 downto 0) := "1110011100011000";
  constant S_BOX_01_43 : std_logic_vector(15 downto 0) := "0010010001111110";
  signal addr_00x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_01_44 : std_logic_vector(15 downto 0) := "0100011110010101";
  constant S_BOX_01_45 : std_logic_vector(15 downto 0) := "0101110100011010";
  constant S_BOX_01_46 : std_logic_vector(15 downto 0) := "1100110000101101";
  constant S_BOX_01_47 : std_logic_vector(15 downto 0) := "1101000111001001";
  -- state 2 and all relevant data to update it
  signal state_02 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #2
  signal addr_01x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_02_00 : std_logic_vector(15 downto 0) := "1101101000000111";
  constant S_BOX_02_01 : std_logic_vector(15 downto 0) := "0010111100010011";
  constant S_BOX_02_02 : std_logic_vector(15 downto 0) := "0110011011000110";
  constant S_BOX_02_03 : std_logic_vector(15 downto 0) := "0111001101001001";
  signal addr_01x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_02_04 : std_logic_vector(15 downto 0) := "1011111011000000";
  constant S_BOX_02_05 : std_logic_vector(15 downto 0) := "1000011101001101";
  constant S_BOX_02_06 : std_logic_vector(15 downto 0) := "1110100001011001";
  constant S_BOX_02_07 : std_logic_vector(15 downto 0) := "1110001010001110";
  signal addr_01x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_02_08 : std_logic_vector(15 downto 0) := "0010111010001011";
  constant S_BOX_02_09 : std_logic_vector(15 downto 0) := "1100111000111000";
  constant S_BOX_02_10 : std_logic_vector(15 downto 0) := "0110010111011000";
  constant S_BOX_02_11 : std_logic_vector(15 downto 0) := "0101011011100001";
  signal addr_01x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_02_12 : std_logic_vector(15 downto 0) := "1000100101110110";
  constant S_BOX_02_13 : std_logic_vector(15 downto 0) := "0101010101100011";
  constant S_BOX_02_14 : std_logic_vector(15 downto 0) := "0011000111010101";
  constant S_BOX_02_15 : std_logic_vector(15 downto 0) := "1011010100001110";
  signal addr_01x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_02_16 : std_logic_vector(15 downto 0) := "1000001101101110";
  constant S_BOX_02_17 : std_logic_vector(15 downto 0) := "0111100101001010";
  constant S_BOX_02_18 : std_logic_vector(15 downto 0) := "1100101110011000";
  constant S_BOX_02_19 : std_logic_vector(15 downto 0) := "1110010011101000";
  signal addr_01x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_02_20 : std_logic_vector(15 downto 0) := "1100101101011000";
  constant S_BOX_02_21 : std_logic_vector(15 downto 0) := "1010001101100101";
  constant S_BOX_02_22 : std_logic_vector(15 downto 0) := "1101111000100100";
  constant S_BOX_02_23 : std_logic_vector(15 downto 0) := "0100011011101001";
  signal addr_01x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_02_24 : std_logic_vector(15 downto 0) := "1100100111100001";
  constant S_BOX_02_25 : std_logic_vector(15 downto 0) := "0110100010010111";
  constant S_BOX_02_26 : std_logic_vector(15 downto 0) := "1100110100001110";
  constant S_BOX_02_27 : std_logic_vector(15 downto 0) := "1001110000110011";
  signal addr_01x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_02_28 : std_logic_vector(15 downto 0) := "1101001100010110";
  constant S_BOX_02_29 : std_logic_vector(15 downto 0) := "1110101000100011";
  constant S_BOX_02_30 : std_logic_vector(15 downto 0) := "1001101010101100";
  constant S_BOX_02_31 : std_logic_vector(15 downto 0) := "0000011110100111";
  signal addr_01x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_02_32 : std_logic_vector(15 downto 0) := "0110100101100011";
  constant S_BOX_02_33 : std_logic_vector(15 downto 0) := "1011011001100010";
  constant S_BOX_02_34 : std_logic_vector(15 downto 0) := "0101010011100101";
  constant S_BOX_02_35 : std_logic_vector(15 downto 0) := "1101000101010110";
  signal addr_01x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_02_36 : std_logic_vector(15 downto 0) := "1010010010111010";
  constant S_BOX_02_37 : std_logic_vector(15 downto 0) := "1110000110001101";
  constant S_BOX_02_38 : std_logic_vector(15 downto 0) := "0110001011110001";
  constant S_BOX_02_39 : std_logic_vector(15 downto 0) := "0100100111011010";
  signal addr_01x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_02_40 : std_logic_vector(15 downto 0) := "1000010111111000";
  constant S_BOX_02_41 : std_logic_vector(15 downto 0) := "0111011001110000";
  constant S_BOX_02_42 : std_logic_vector(15 downto 0) := "0011110101001100";
  constant S_BOX_02_43 : std_logic_vector(15 downto 0) := "0101000011101101";
  signal addr_01x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_02_44 : std_logic_vector(15 downto 0) := "0101010101110100";
  constant S_BOX_02_45 : std_logic_vector(15 downto 0) := "0101101001010011";
  constant S_BOX_02_46 : std_logic_vector(15 downto 0) := "1000011011110010";
  constant S_BOX_02_47 : std_logic_vector(15 downto 0) := "1001000000111111";
  -- state 3 and all relevant data to update it
  signal state_03 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #3
  signal addr_02x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_03_00 : std_logic_vector(15 downto 0) := "0101000111001011";
  constant S_BOX_03_01 : std_logic_vector(15 downto 0) := "0110000101110101";
  constant S_BOX_03_02 : std_logic_vector(15 downto 0) := "1101100100010110";
  constant S_BOX_03_03 : std_logic_vector(15 downto 0) := "0001110110100101";
  signal addr_02x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_03_04 : std_logic_vector(15 downto 0) := "0011010110000111";
  constant S_BOX_03_05 : std_logic_vector(15 downto 0) := "1000000011110111";
  constant S_BOX_03_06 : std_logic_vector(15 downto 0) := "0101110001010101";
  constant S_BOX_03_07 : std_logic_vector(15 downto 0) := "0011101011100100";
  signal addr_02x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_03_08 : std_logic_vector(15 downto 0) := "1001111000001011";
  constant S_BOX_03_09 : std_logic_vector(15 downto 0) := "1010011101010010";
  constant S_BOX_03_10 : std_logic_vector(15 downto 0) := "0111011100100001";
  constant S_BOX_03_11 : std_logic_vector(15 downto 0) := "0110010010011011";
  signal addr_02x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_03_12 : std_logic_vector(15 downto 0) := "1001010111110000";
  constant S_BOX_03_13 : std_logic_vector(15 downto 0) := "0010010101011011";
  constant S_BOX_03_14 : std_logic_vector(15 downto 0) := "0010001110110101";
  constant S_BOX_03_15 : std_logic_vector(15 downto 0) := "0111000101100110";
  signal addr_02x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_03_16 : std_logic_vector(15 downto 0) := "1100111000011001";
  constant S_BOX_03_17 : std_logic_vector(15 downto 0) := "0110011100001110";
  constant S_BOX_03_18 : std_logic_vector(15 downto 0) := "1000011111010010";
  constant S_BOX_03_19 : std_logic_vector(15 downto 0) := "0011110110011000";
  signal addr_02x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_03_20 : std_logic_vector(15 downto 0) := "0001100111111000";
  constant S_BOX_03_21 : std_logic_vector(15 downto 0) := "0010101010110101";
  constant S_BOX_03_22 : std_logic_vector(15 downto 0) := "1000111100101001";
  constant S_BOX_03_23 : std_logic_vector(15 downto 0) := "1111100000011001";
  signal addr_02x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_03_24 : std_logic_vector(15 downto 0) := "1001111100100001";
  constant S_BOX_03_25 : std_logic_vector(15 downto 0) := "1011010000111100";
  constant S_BOX_03_26 : std_logic_vector(15 downto 0) := "0100011000101111";
  constant S_BOX_03_27 : std_logic_vector(15 downto 0) := "0101111001010100";
  signal addr_02x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_03_28 : std_logic_vector(15 downto 0) := "0011101010010011";
  constant S_BOX_03_29 : std_logic_vector(15 downto 0) := "1110010000010111";
  constant S_BOX_03_30 : std_logic_vector(15 downto 0) := "0110110110100001";
  constant S_BOX_03_31 : std_logic_vector(15 downto 0) := "0111100100011100";
  signal addr_02x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_03_32 : std_logic_vector(15 downto 0) := "0000101110101110";
  constant S_BOX_03_33 : std_logic_vector(15 downto 0) := "1100011011101000";
  constant S_BOX_03_34 : std_logic_vector(15 downto 0) := "0001110001101101";
  constant S_BOX_03_35 : std_logic_vector(15 downto 0) := "0100100111011001";
  signal addr_02x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_03_36 : std_logic_vector(15 downto 0) := "1000011111011000";
  constant S_BOX_03_37 : std_logic_vector(15 downto 0) := "0110001001011110";
  constant S_BOX_03_38 : std_logic_vector(15 downto 0) := "0101011010010101";
  constant S_BOX_03_39 : std_logic_vector(15 downto 0) := "1000110001010111";
  signal addr_02x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_03_40 : std_logic_vector(15 downto 0) := "1001110000011011";
  constant S_BOX_03_41 : std_logic_vector(15 downto 0) := "1010011001110001";
  constant S_BOX_03_42 : std_logic_vector(15 downto 0) := "1000111110100010";
  constant S_BOX_03_43 : std_logic_vector(15 downto 0) := "1111101010010000";
  signal addr_02x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_03_44 : std_logic_vector(15 downto 0) := "0001110010011110";
  constant S_BOX_03_45 : std_logic_vector(15 downto 0) := "1111110000100100";
  constant S_BOX_03_46 : std_logic_vector(15 downto 0) := "1000110100101011";
  constant S_BOX_03_47 : std_logic_vector(15 downto 0) := "0101011100110010";
  -- state 4 and all relevant data to update it
  signal state_04 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #4
  signal addr_03x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_04_00 : std_logic_vector(15 downto 0) := "0110011001011100";
  constant S_BOX_04_01 : std_logic_vector(15 downto 0) := "1110010100101010";
  constant S_BOX_04_02 : std_logic_vector(15 downto 0) := "0011000111101100";
  constant S_BOX_04_03 : std_logic_vector(15 downto 0) := "1010010010110101";
  signal addr_03x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_04_04 : std_logic_vector(15 downto 0) := "1010111000101100";
  constant S_BOX_04_05 : std_logic_vector(15 downto 0) := "1100001011011100";
  constant S_BOX_04_06 : std_logic_vector(15 downto 0) := "1000110111001010";
  constant S_BOX_04_07 : std_logic_vector(15 downto 0) := "1100100010100111";
  signal addr_03x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_04_08 : std_logic_vector(15 downto 0) := "0110101010001101";
  constant S_BOX_04_09 : std_logic_vector(15 downto 0) := "0011001100100111";
  constant S_BOX_04_10 : std_logic_vector(15 downto 0) := "1011101100011000";
  constant S_BOX_04_11 : std_logic_vector(15 downto 0) := "0100111100010011";
  signal addr_03x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_04_12 : std_logic_vector(15 downto 0) := "0101110001110100";
  constant S_BOX_04_13 : std_logic_vector(15 downto 0) := "1111100010000110";
  constant S_BOX_04_14 : std_logic_vector(15 downto 0) := "0000110010101111";
  constant S_BOX_04_15 : std_logic_vector(15 downto 0) := "1001101001100011";
  signal addr_03x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_04_16 : std_logic_vector(15 downto 0) := "1001011100110001";
  constant S_BOX_04_17 : std_logic_vector(15 downto 0) := "1111010001000101";
  constant S_BOX_04_18 : std_logic_vector(15 downto 0) := "0101011101001010";
  constant S_BOX_04_19 : std_logic_vector(15 downto 0) := "0110110100100011";
  signal addr_03x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_04_20 : std_logic_vector(15 downto 0) := "1010101001001110";
  constant S_BOX_04_21 : std_logic_vector(15 downto 0) := "0100110001111010";
  constant S_BOX_04_22 : std_logic_vector(15 downto 0) := "0110000101100111";
  constant S_BOX_04_23 : std_logic_vector(15 downto 0) := "1111100000010011";
  signal addr_03x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_04_24 : std_logic_vector(15 downto 0) := "0110001001101011";
  constant S_BOX_04_25 : std_logic_vector(15 downto 0) := "0000011111101100";
  constant S_BOX_04_26 : std_logic_vector(15 downto 0) := "1000011011010011";
  constant S_BOX_04_27 : std_logic_vector(15 downto 0) := "1010111000001110";
  signal addr_03x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_04_28 : std_logic_vector(15 downto 0) := "1110100100001101";
  constant S_BOX_04_29 : std_logic_vector(15 downto 0) := "1010011101000011";
  constant S_BOX_04_30 : std_logic_vector(15 downto 0) := "0000110111011001";
  constant S_BOX_04_31 : std_logic_vector(15 downto 0) := "0010011000111101";
  signal addr_03x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_04_32 : std_logic_vector(15 downto 0) := "0111010010010110";
  constant S_BOX_04_33 : std_logic_vector(15 downto 0) := "0011110101001010";
  constant S_BOX_04_34 : std_logic_vector(15 downto 0) := "1110011100001100";
  constant S_BOX_04_35 : std_logic_vector(15 downto 0) := "1111100110000001";
  signal addr_03x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_04_36 : std_logic_vector(15 downto 0) := "1010101110000011";
  constant S_BOX_04_37 : std_logic_vector(15 downto 0) := "0011111100101000";
  constant S_BOX_04_38 : std_logic_vector(15 downto 0) := "0001001110011101";
  constant S_BOX_04_39 : std_logic_vector(15 downto 0) := "0111001000100111";
  signal addr_03x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_04_40 : std_logic_vector(15 downto 0) := "0010100100111011";
  constant S_BOX_04_41 : std_logic_vector(15 downto 0) := "1011010010010011";
  constant S_BOX_04_42 : std_logic_vector(15 downto 0) := "0011011101001010";
  constant S_BOX_04_43 : std_logic_vector(15 downto 0) := "0011000011101101";
  signal addr_03x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_04_44 : std_logic_vector(15 downto 0) := "0100110101010101";
  constant S_BOX_04_45 : std_logic_vector(15 downto 0) := "1000010011111001";
  constant S_BOX_04_46 : std_logic_vector(15 downto 0) := "1111000101011000";
  constant S_BOX_04_47 : std_logic_vector(15 downto 0) := "1001111111000000";
  -- state 5 and all relevant data to update it
  signal state_05 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #5
  signal addr_04x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_05_00 : std_logic_vector(15 downto 0) := "1101111000100010";
  constant S_BOX_05_01 : std_logic_vector(15 downto 0) := "0010111110000110";
  constant S_BOX_05_02 : std_logic_vector(15 downto 0) := "1011110000011100";
  constant S_BOX_05_03 : std_logic_vector(15 downto 0) := "0001100101110110";
  signal addr_04x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_05_04 : std_logic_vector(15 downto 0) := "0011010010111001";
  constant S_BOX_05_05 : std_logic_vector(15 downto 0) := "0100110011011100";
  constant S_BOX_05_06 : std_logic_vector(15 downto 0) := "1000010101110101";
  constant S_BOX_05_07 : std_logic_vector(15 downto 0) := "1101011011100000";
  signal addr_04x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_05_08 : std_logic_vector(15 downto 0) := "1110100000011011";
  constant S_BOX_05_09 : std_logic_vector(15 downto 0) := "1111011000000101";
  constant S_BOX_05_10 : std_logic_vector(15 downto 0) := "0101101001110001";
  constant S_BOX_05_11 : std_logic_vector(15 downto 0) := "1001010100110011";
  signal addr_04x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_05_12 : std_logic_vector(15 downto 0) := "0110111001000101";
  constant S_BOX_05_13 : std_logic_vector(15 downto 0) := "0001110011011001";
  constant S_BOX_05_14 : std_logic_vector(15 downto 0) := "1010011010101001";
  constant S_BOX_05_15 : std_logic_vector(15 downto 0) := "1100001111010001";
  signal addr_04x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_05_16 : std_logic_vector(15 downto 0) := "1010111010000101";
  constant S_BOX_05_17 : std_logic_vector(15 downto 0) := "1100110110101000";
  constant S_BOX_05_18 : std_logic_vector(15 downto 0) := "0011100111100001";
  constant S_BOX_05_19 : std_logic_vector(15 downto 0) := "0101110000100111";
  signal addr_04x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_05_20 : std_logic_vector(15 downto 0) := "1100010101100011";
  constant S_BOX_05_21 : std_logic_vector(15 downto 0) := "0010011100010111";
  constant S_BOX_05_22 : std_logic_vector(15 downto 0) := "1010100001011011";
  constant S_BOX_05_23 : std_logic_vector(15 downto 0) := "0111111001000001";
  signal addr_04x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_05_24 : std_logic_vector(15 downto 0) := "1001011110011000";
  constant S_BOX_05_25 : std_logic_vector(15 downto 0) := "1010110110100001";
  constant S_BOX_05_26 : std_logic_vector(15 downto 0) := "1001100011101100";
  constant S_BOX_05_27 : std_logic_vector(15 downto 0) := "1110101100001100";
  signal addr_04x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_05_28 : std_logic_vector(15 downto 0) := "1100011010011001";
  constant S_BOX_05_29 : std_logic_vector(15 downto 0) := "0101001111001010";
  constant S_BOX_05_30 : std_logic_vector(15 downto 0) := "0100111001100011";
  constant S_BOX_05_31 : std_logic_vector(15 downto 0) := "1011101001001001";
  signal addr_04x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_05_32 : std_logic_vector(15 downto 0) := "1111011110000000";
  constant S_BOX_05_33 : std_logic_vector(15 downto 0) := "1010100110100011";
  constant S_BOX_05_34 : std_logic_vector(15 downto 0) := "0011110010011010";
  constant S_BOX_05_35 : std_logic_vector(15 downto 0) := "0010011100010111";
  signal addr_04x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_05_36 : std_logic_vector(15 downto 0) := "1100111001010001";
  constant S_BOX_05_37 : std_logic_vector(15 downto 0) := "0010111000111100";
  constant S_BOX_05_38 : std_logic_vector(15 downto 0) := "0100001110011101";
  constant S_BOX_05_39 : std_logic_vector(15 downto 0) := "0101100011110100";
  signal addr_04x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_05_40 : std_logic_vector(15 downto 0) := "1000110010001111";
  constant S_BOX_05_41 : std_logic_vector(15 downto 0) := "0100011011010011";
  constant S_BOX_05_42 : std_logic_vector(15 downto 0) := "0110100000110111";
  constant S_BOX_05_43 : std_logic_vector(15 downto 0) := "1001001010110110";
  signal addr_04x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_05_44 : std_logic_vector(15 downto 0) := "0001100001111110";
  constant S_BOX_05_45 : std_logic_vector(15 downto 0) := "0010111011010100";
  constant S_BOX_05_46 : std_logic_vector(15 downto 0) := "1110110000100110";
  constant S_BOX_05_47 : std_logic_vector(15 downto 0) := "1011000111000110";
  -- state 6 and all relevant data to update it
  signal state_06 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #6
  signal addr_05x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_06_00 : std_logic_vector(15 downto 0) := "1101000101101100";
  constant S_BOX_06_01 : std_logic_vector(15 downto 0) := "1111010011010000";
  constant S_BOX_06_02 : std_logic_vector(15 downto 0) := "1011100000111010";
  constant S_BOX_06_03 : std_logic_vector(15 downto 0) := "1110110000001101";
  signal addr_05x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_06_04 : std_logic_vector(15 downto 0) := "0001011000011111";
  constant S_BOX_06_05 : std_logic_vector(15 downto 0) := "1011110100011000";
  constant S_BOX_06_06 : std_logic_vector(15 downto 0) := "1000110001110101";
  constant S_BOX_06_07 : std_logic_vector(15 downto 0) := "1110011001001001";
  signal addr_05x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_06_08 : std_logic_vector(15 downto 0) := "1000111000111100";
  constant S_BOX_06_09 : std_logic_vector(15 downto 0) := "0011110101100100";
  constant S_BOX_06_10 : std_logic_vector(15 downto 0) := "1101000110101100";
  constant S_BOX_06_11 : std_logic_vector(15 downto 0) := "0010010110111010";
  signal addr_05x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_06_12 : std_logic_vector(15 downto 0) := "0110011100010110";
  constant S_BOX_06_13 : std_logic_vector(15 downto 0) := "0000001001111111";
  constant S_BOX_06_14 : std_logic_vector(15 downto 0) := "1011011000001011";
  constant S_BOX_06_15 : std_logic_vector(15 downto 0) := "1000011111010001";
  signal addr_05x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_06_16 : std_logic_vector(15 downto 0) := "1111100000101001";
  constant S_BOX_06_17 : std_logic_vector(15 downto 0) := "1100101111001000";
  constant S_BOX_06_18 : std_logic_vector(15 downto 0) := "1101010011010001";
  constant S_BOX_06_19 : std_logic_vector(15 downto 0) := "1010001001011011";
  signal addr_05x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_06_20 : std_logic_vector(15 downto 0) := "0110101001100110";
  constant S_BOX_06_21 : std_logic_vector(15 downto 0) := "1110000101010011";
  constant S_BOX_06_22 : std_logic_vector(15 downto 0) := "1101101001001001";
  constant S_BOX_06_23 : std_logic_vector(15 downto 0) := "1010011001011100";
  signal addr_05x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_06_24 : std_logic_vector(15 downto 0) := "1111110010010000";
  constant S_BOX_06_25 : std_logic_vector(15 downto 0) := "0111010001000111";
  constant S_BOX_06_26 : std_logic_vector(15 downto 0) := "0011001011011001";
  constant S_BOX_06_27 : std_logic_vector(15 downto 0) := "1010011101010010";
  signal addr_05x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_06_28 : std_logic_vector(15 downto 0) := "1010101010001101";
  constant S_BOX_06_29 : std_logic_vector(15 downto 0) := "1110001011010010";
  constant S_BOX_06_30 : std_logic_vector(15 downto 0) := "1010010000110111";
  constant S_BOX_06_31 : std_logic_vector(15 downto 0) := "1001100011100011";
  signal addr_05x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_06_32 : std_logic_vector(15 downto 0) := "0011011010101010";
  constant S_BOX_06_33 : std_logic_vector(15 downto 0) := "1101000000111011";
  constant S_BOX_06_34 : std_logic_vector(15 downto 0) := "1001101010011100";
  constant S_BOX_06_35 : std_logic_vector(15 downto 0) := "1001011100100101";
  signal addr_05x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_06_36 : std_logic_vector(15 downto 0) := "0010111101001001";
  constant S_BOX_06_37 : std_logic_vector(15 downto 0) := "1101101100010001";
  constant S_BOX_06_38 : std_logic_vector(15 downto 0) := "1010011000010111";
  constant S_BOX_06_39 : std_logic_vector(15 downto 0) := "0001010111010011";
  signal addr_05x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_06_40 : std_logic_vector(15 downto 0) := "0101000101110011";
  constant S_BOX_06_41 : std_logic_vector(15 downto 0) := "1111001010100010";
  constant S_BOX_06_42 : std_logic_vector(15 downto 0) := "1101100011001001";
  constant S_BOX_06_43 : std_logic_vector(15 downto 0) := "0100111110100001";
  signal addr_05x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_06_44 : std_logic_vector(15 downto 0) := "1000011101100011";
  constant S_BOX_06_45 : std_logic_vector(15 downto 0) := "0100100101110110";
  constant S_BOX_06_46 : std_logic_vector(15 downto 0) := "0010111001001110";
  constant S_BOX_06_47 : std_logic_vector(15 downto 0) := "1110110010100010";
  -- state 7 and all relevant data to update it
  signal state_07 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #7
  signal addr_06x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_07_00 : std_logic_vector(15 downto 0) := "0100011111001010";
  constant S_BOX_07_01 : std_logic_vector(15 downto 0) := "1110010000001111";
  constant S_BOX_07_02 : std_logic_vector(15 downto 0) := "1010110011010010";
  constant S_BOX_07_03 : std_logic_vector(15 downto 0) := "1101011010010100";
  signal addr_06x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_07_04 : std_logic_vector(15 downto 0) := "0000010110111011";
  constant S_BOX_07_05 : std_logic_vector(15 downto 0) := "0110101100001011";
  constant S_BOX_07_06 : std_logic_vector(15 downto 0) := "1011110010001010";
  constant S_BOX_07_07 : std_logic_vector(15 downto 0) := "0011001011010011";
  signal addr_06x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_07_08 : std_logic_vector(15 downto 0) := "0110011111000010";
  constant S_BOX_07_09 : std_logic_vector(15 downto 0) := "0110100101101100";
  constant S_BOX_07_10 : std_logic_vector(15 downto 0) := "1011010011001100";
  constant S_BOX_07_11 : std_logic_vector(15 downto 0) := "1110110000011010";
  signal addr_06x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_07_12 : std_logic_vector(15 downto 0) := "1001110100110100";
  constant S_BOX_07_13 : std_logic_vector(15 downto 0) := "1100100010010111";
  constant S_BOX_07_14 : std_logic_vector(15 downto 0) := "1011000010101101";
  constant S_BOX_07_15 : std_logic_vector(15 downto 0) := "1101110001001001";
  signal addr_06x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_07_16 : std_logic_vector(15 downto 0) := "0101011100011100";
  constant S_BOX_07_17 : std_logic_vector(15 downto 0) := "1100001011110100";
  constant S_BOX_07_18 : std_logic_vector(15 downto 0) := "1101110000110001";
  constant S_BOX_07_19 : std_logic_vector(15 downto 0) := "0100110001101110";
  signal addr_06x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_07_20 : std_logic_vector(15 downto 0) := "1110010100101001";
  constant S_BOX_07_21 : std_logic_vector(15 downto 0) := "0001100111101001";
  constant S_BOX_07_22 : std_logic_vector(15 downto 0) := "1000110001011011";
  constant S_BOX_07_23 : std_logic_vector(15 downto 0) := "0011011101010001";
  signal addr_06x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_07_24 : std_logic_vector(15 downto 0) := "0001110111001001";
  constant S_BOX_07_25 : std_logic_vector(15 downto 0) := "1000101101010011";
  constant S_BOX_07_26 : std_logic_vector(15 downto 0) := "1000011111100100";
  constant S_BOX_07_27 : std_logic_vector(15 downto 0) := "0010111100001110";
  signal addr_06x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_07_28 : std_logic_vector(15 downto 0) := "1100000101111001";
  constant S_BOX_07_29 : std_logic_vector(15 downto 0) := "1010101001110010";
  constant S_BOX_07_30 : std_logic_vector(15 downto 0) := "1000111001001101";
  constant S_BOX_07_31 : std_logic_vector(15 downto 0) := "0001011101011010";
  signal addr_06x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_07_32 : std_logic_vector(15 downto 0) := "0011101010110010";
  constant S_BOX_07_33 : std_logic_vector(15 downto 0) := "0101010010110101";
  constant S_BOX_07_34 : std_logic_vector(15 downto 0) := "0011000100101111";
  constant S_BOX_07_35 : std_logic_vector(15 downto 0) := "1110001100110100";
  signal addr_06x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_07_36 : std_logic_vector(15 downto 0) := "1011101000001101";
  constant S_BOX_07_37 : std_logic_vector(15 downto 0) := "0010110010110101";
  constant S_BOX_07_38 : std_logic_vector(15 downto 0) := "0101101110010001";
  constant S_BOX_07_39 : std_logic_vector(15 downto 0) := "1010101100110010";
  signal addr_06x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_07_40 : std_logic_vector(15 downto 0) := "1000010100111101";
  constant S_BOX_07_41 : std_logic_vector(15 downto 0) := "0101110000011110";
  constant S_BOX_07_42 : std_logic_vector(15 downto 0) := "0010111100000111";
  constant S_BOX_07_43 : std_logic_vector(15 downto 0) := "0011010101101010";
  signal addr_06x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_07_44 : std_logic_vector(15 downto 0) := "1001110100110100";
  constant S_BOX_07_45 : std_logic_vector(15 downto 0) := "0011000101111001";
  constant S_BOX_07_46 : std_logic_vector(15 downto 0) := "1010101100010011";
  constant S_BOX_07_47 : std_logic_vector(15 downto 0) := "1000011111100001";
  -- state 8 and all relevant data to update it
  signal state_08 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #8
  signal addr_07x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_08_00 : std_logic_vector(15 downto 0) := "0110111011000001";
  constant S_BOX_08_01 : std_logic_vector(15 downto 0) := "0010001101010111";
  constant S_BOX_08_02 : std_logic_vector(15 downto 0) := "1111000110000011";
  constant S_BOX_08_03 : std_logic_vector(15 downto 0) := "1100101100011001";
  signal addr_07x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_08_04 : std_logic_vector(15 downto 0) := "1101000111100100";
  constant S_BOX_08_05 : std_logic_vector(15 downto 0) := "1010011111000001";
  constant S_BOX_08_06 : std_logic_vector(15 downto 0) := "0101010011001011";
  constant S_BOX_08_07 : std_logic_vector(15 downto 0) := "1011010001111000";
  signal addr_07x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_08_08 : std_logic_vector(15 downto 0) := "1110110101010000";
  constant S_BOX_08_09 : std_logic_vector(15 downto 0) := "0101010110011010";
  constant S_BOX_08_10 : std_logic_vector(15 downto 0) := "1000110000011111";
  constant S_BOX_08_11 : std_logic_vector(15 downto 0) := "1111010000101001";
  signal addr_07x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_08_12 : std_logic_vector(15 downto 0) := "0111111100001000";
  constant S_BOX_08_13 : std_logic_vector(15 downto 0) := "0011001011011001";
  constant S_BOX_08_14 : std_logic_vector(15 downto 0) := "1010100110001011";
  constant S_BOX_08_15 : std_logic_vector(15 downto 0) := "0010011100010111";
  signal addr_07x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_08_16 : std_logic_vector(15 downto 0) := "0110001000111101";
  constant S_BOX_08_17 : std_logic_vector(15 downto 0) := "0000011111011001";
  constant S_BOX_08_18 : std_logic_vector(15 downto 0) := "0011101101010100";
  constant S_BOX_08_19 : std_logic_vector(15 downto 0) := "1010110100110001";
  signal addr_07x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_08_20 : std_logic_vector(15 downto 0) := "0110001110110001";
  constant S_BOX_08_21 : std_logic_vector(15 downto 0) := "0001111010100101";
  constant S_BOX_08_22 : std_logic_vector(15 downto 0) := "0110110001101001";
  constant S_BOX_08_23 : std_logic_vector(15 downto 0) := "1101101100001001";
  signal addr_07x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_08_24 : std_logic_vector(15 downto 0) := "0011001110111000";
  constant S_BOX_08_25 : std_logic_vector(15 downto 0) := "1110001010010110";
  constant S_BOX_08_26 : std_logic_vector(15 downto 0) := "0000111010101110";
  constant S_BOX_08_27 : std_logic_vector(15 downto 0) := "0100011101110100";
  signal addr_07x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_08_28 : std_logic_vector(15 downto 0) := "0011010101000111";
  constant S_BOX_08_29 : std_logic_vector(15 downto 0) := "0010001001111101";
  constant S_BOX_08_30 : std_logic_vector(15 downto 0) := "1010011010001110";
  constant S_BOX_08_31 : std_logic_vector(15 downto 0) := "1101000000011111";
  signal addr_07x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_08_32 : std_logic_vector(15 downto 0) := "1011110000011100";
  constant S_BOX_08_33 : std_logic_vector(15 downto 0) := "1110010101110000";
  constant S_BOX_08_34 : std_logic_vector(15 downto 0) := "1100101100011010";
  constant S_BOX_08_35 : std_logic_vector(15 downto 0) := "0101011000111001";
  signal addr_07x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_08_36 : std_logic_vector(15 downto 0) := "1011001011010001";
  constant S_BOX_08_37 : std_logic_vector(15 downto 0) := "0011101110000110";
  constant S_BOX_08_38 : std_logic_vector(15 downto 0) := "1111100000100011";
  constant S_BOX_08_39 : std_logic_vector(15 downto 0) := "0101001101001011";
  signal addr_07x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_08_40 : std_logic_vector(15 downto 0) := "0001011010110011";
  constant S_BOX_08_41 : std_logic_vector(15 downto 0) := "1010010001101011";
  constant S_BOX_08_42 : std_logic_vector(15 downto 0) := "0111011100001010";
  constant S_BOX_08_43 : std_logic_vector(15 downto 0) := "0111000001010111";
  signal addr_07x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_08_44 : std_logic_vector(15 downto 0) := "0100110001100111";
  constant S_BOX_08_45 : std_logic_vector(15 downto 0) := "0001011011101010";
  constant S_BOX_08_46 : std_logic_vector(15 downto 0) := "0011001000110111";
  constant S_BOX_08_47 : std_logic_vector(15 downto 0) := "1100011000111001";
  -- state 9 and all relevant data to update it
  signal state_09 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #9
  signal addr_08x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_09_00 : std_logic_vector(15 downto 0) := "0111001011010010";
  constant S_BOX_09_01 : std_logic_vector(15 downto 0) := "1111010010100001";
  constant S_BOX_09_02 : std_logic_vector(15 downto 0) := "0100110010110110";
  constant S_BOX_09_03 : std_logic_vector(15 downto 0) := "1010101010111000";
  signal addr_08x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_09_04 : std_logic_vector(15 downto 0) := "0111100000011011";
  constant S_BOX_09_05 : std_logic_vector(15 downto 0) := "0011011101001010";
  constant S_BOX_09_06 : std_logic_vector(15 downto 0) := "1000101110011010";
  constant S_BOX_09_07 : std_logic_vector(15 downto 0) := "1010001001110011";
  signal addr_08x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_09_08 : std_logic_vector(15 downto 0) := "0000111001011011";
  constant S_BOX_09_09 : std_logic_vector(15 downto 0) := "1110101001001100";
  constant S_BOX_09_10 : std_logic_vector(15 downto 0) := "0011001100011101";
  constant S_BOX_09_11 : std_logic_vector(15 downto 0) := "0111011001110000";
  signal addr_08x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_09_12 : std_logic_vector(15 downto 0) := "0011010001011011";
  constant S_BOX_09_13 : std_logic_vector(15 downto 0) := "0110001101010110";
  constant S_BOX_09_14 : std_logic_vector(15 downto 0) := "1100010101101010";
  constant S_BOX_09_15 : std_logic_vector(15 downto 0) := "0001000111111100";
  signal addr_08x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_09_16 : std_logic_vector(15 downto 0) := "0010111011000011";
  constant S_BOX_09_17 : std_logic_vector(15 downto 0) := "1001111010001100";
  constant S_BOX_09_18 : std_logic_vector(15 downto 0) := "1001001110100011";
  constant S_BOX_09_19 : std_logic_vector(15 downto 0) := "0001101001110101";
  signal addr_08x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_09_20 : std_logic_vector(15 downto 0) := "0000100011111011";
  constant S_BOX_09_21 : std_logic_vector(15 downto 0) := "1110000111011000";
  constant S_BOX_09_22 : std_logic_vector(15 downto 0) := "1010010001010111";
  constant S_BOX_09_23 : std_logic_vector(15 downto 0) := "0011100110010101";
  signal addr_08x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_09_24 : std_logic_vector(15 downto 0) := "0010011110011001";
  constant S_BOX_09_25 : std_logic_vector(15 downto 0) := "0110100100111100";
  constant S_BOX_09_26 : std_logic_vector(15 downto 0) := "1100001011011100";
  constant S_BOX_09_27 : std_logic_vector(15 downto 0) := "0001000111110101";
  signal addr_08x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_09_28 : std_logic_vector(15 downto 0) := "0110100110100101";
  constant S_BOX_09_29 : std_logic_vector(15 downto 0) := "1100001101010101";
  constant S_BOX_09_30 : std_logic_vector(15 downto 0) := "1101100100111000";
  constant S_BOX_09_31 : std_logic_vector(15 downto 0) := "0011010101110001";
  signal addr_08x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_09_32 : std_logic_vector(15 downto 0) := "1000101111101000";
  constant S_BOX_09_33 : std_logic_vector(15 downto 0) := "1011000011110100";
  constant S_BOX_09_34 : std_logic_vector(15 downto 0) := "0010001111010011";
  constant S_BOX_09_35 : std_logic_vector(15 downto 0) := "0110101001100110";
  signal addr_08x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_09_36 : std_logic_vector(15 downto 0) := "0110110110001001";
  constant S_BOX_09_37 : std_logic_vector(15 downto 0) := "0100100011110011";
  constant S_BOX_09_38 : std_logic_vector(15 downto 0) := "1101110001011000";
  constant S_BOX_09_39 : std_logic_vector(15 downto 0) := "0011101000111001";
  signal addr_08x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_09_40 : std_logic_vector(15 downto 0) := "0011001011101100";
  constant S_BOX_09_41 : std_logic_vector(15 downto 0) := "0011100101010110";
  constant S_BOX_09_42 : std_logic_vector(15 downto 0) := "1110101101100000";
  constant S_BOX_09_43 : std_logic_vector(15 downto 0) := "0101011111000010";
  signal addr_08x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_09_44 : std_logic_vector(15 downto 0) := "0010001001111101";
  constant S_BOX_09_45 : std_logic_vector(15 downto 0) := "1100011000010111";
  constant S_BOX_09_46 : std_logic_vector(15 downto 0) := "0110111010011000";
  constant S_BOX_09_47 : std_logic_vector(15 downto 0) := "1000111101001001";
  -- state 10 and all relevant data to update it
  signal state_10 : std_logic_vector(47 downto 0) := SEED; -- scrambling stage #10
  signal addr_09x_00 : std_logic_vector(3 downto 0);
  constant S_BOX_10_00 : std_logic_vector(15 downto 0) := "0000111011100110";
  constant S_BOX_10_01 : std_logic_vector(15 downto 0) := "1101010111000100";
  constant S_BOX_10_02 : std_logic_vector(15 downto 0) := "0101111000010101";
  constant S_BOX_10_03 : std_logic_vector(15 downto 0) := "0001011110011010";
  signal addr_09x_01 : std_logic_vector(3 downto 0);
  constant S_BOX_10_04 : std_logic_vector(15 downto 0) := "1010010100101011";
  constant S_BOX_10_05 : std_logic_vector(15 downto 0) := "0111100100001101";
  constant S_BOX_10_06 : std_logic_vector(15 downto 0) := "0001011000111101";
  constant S_BOX_10_07 : std_logic_vector(15 downto 0) := "1100001110100101";
  signal addr_09x_02 : std_logic_vector(3 downto 0);
  constant S_BOX_10_08 : std_logic_vector(15 downto 0) := "0101011001110100";
  constant S_BOX_10_09 : std_logic_vector(15 downto 0) := "1100100001110011";
  constant S_BOX_10_10 : std_logic_vector(15 downto 0) := "1100010110010101";
  constant S_BOX_10_11 : std_logic_vector(15 downto 0) := "1100101100101100";
  signal addr_09x_03 : std_logic_vector(3 downto 0);
  constant S_BOX_10_12 : std_logic_vector(15 downto 0) := "1110001001110001";
  constant S_BOX_10_13 : std_logic_vector(15 downto 0) := "1101011100000011";
  constant S_BOX_10_14 : std_logic_vector(15 downto 0) := "1010011010101010";
  constant S_BOX_10_15 : std_logic_vector(15 downto 0) := "0011011011000101";
  signal addr_09x_04 : std_logic_vector(3 downto 0);
  constant S_BOX_10_16 : std_logic_vector(15 downto 0) := "1000000011111101";
  constant S_BOX_10_17 : std_logic_vector(15 downto 0) := "1011101001010001";
  constant S_BOX_10_18 : std_logic_vector(15 downto 0) := "1010011101001100";
  constant S_BOX_10_19 : std_logic_vector(15 downto 0) := "0101001101100101";
  signal addr_09x_05 : std_logic_vector(3 downto 0);
  constant S_BOX_10_20 : std_logic_vector(15 downto 0) := "0010111110000110";
  constant S_BOX_10_21 : std_logic_vector(15 downto 0) := "0100100110111010";
  constant S_BOX_10_22 : std_logic_vector(15 downto 0) := "1111001110010000";
  constant S_BOX_10_23 : std_logic_vector(15 downto 0) := "0001101010110101";
  signal addr_09x_06 : std_logic_vector(3 downto 0);
  constant S_BOX_10_24 : std_logic_vector(15 downto 0) := "1100010000111011";
  constant S_BOX_10_25 : std_logic_vector(15 downto 0) := "0000110101111100";
  constant S_BOX_10_26 : std_logic_vector(15 downto 0) := "0101001100011110";
  constant S_BOX_10_27 : std_logic_vector(15 downto 0) := "1001000111110010";
  signal addr_09x_07 : std_logic_vector(3 downto 0);
  constant S_BOX_10_28 : std_logic_vector(15 downto 0) := "0001000111010111";
  constant S_BOX_10_29 : std_logic_vector(15 downto 0) := "0011011000011110";
  constant S_BOX_10_30 : std_logic_vector(15 downto 0) := "0011110001100011";
  constant S_BOX_10_31 : std_logic_vector(15 downto 0) := "1000111010010011";
  signal addr_09x_08 : std_logic_vector(3 downto 0);
  constant S_BOX_10_32 : std_logic_vector(15 downto 0) := "0011001110111000";
  constant S_BOX_10_33 : std_logic_vector(15 downto 0) := "0101111111000000";
  constant S_BOX_10_34 : std_logic_vector(15 downto 0) := "1101011000011001";
  constant S_BOX_10_35 : std_logic_vector(15 downto 0) := "0011010011010011";
  signal addr_09x_09 : std_logic_vector(3 downto 0);
  constant S_BOX_10_36 : std_logic_vector(15 downto 0) := "0111010010100110";
  constant S_BOX_10_37 : std_logic_vector(15 downto 0) := "0011110000011101";
  constant S_BOX_10_38 : std_logic_vector(15 downto 0) := "1111100001110000";
  constant S_BOX_10_39 : std_logic_vector(15 downto 0) := "0101011001010011";
  signal addr_09x_10 : std_logic_vector(3 downto 0);
  constant S_BOX_10_40 : std_logic_vector(15 downto 0) := "1100101110001010";
  constant S_BOX_10_41 : std_logic_vector(15 downto 0) := "1001010100111010";
  constant S_BOX_10_42 : std_logic_vector(15 downto 0) := "1011101000100110";
  constant S_BOX_10_43 : std_logic_vector(15 downto 0) := "0010100011111010";
  signal addr_09x_11 : std_logic_vector(3 downto 0);
  constant S_BOX_10_44 : std_logic_vector(15 downto 0) := "0111111000001010";
  constant S_BOX_10_45 : std_logic_vector(15 downto 0) := "0010011001111001";
  constant S_BOX_10_46 : std_logic_vector(15 downto 0) := "1110100101001001";
  constant S_BOX_10_47 : std_logic_vector(15 downto 0) := "0100010110011011";
begin
  --
  -- Output
  --
  rnd <= state_10(N_BITS-1 downto 0); -- warning: do not use in the very first 10 clock cycles (not random enough)
  --
  -- S-box addresses (P-boxes)
  --
  addr_00x_00 <= state_00(24) & state_00(40) & state_00(41) & state_00(26);
  addr_00x_01 <= state_00( 7) & state_00(10) & state_00(15) & state_00(36);
  addr_00x_02 <= state_00(34) & state_00(32) & state_00(38) & state_00(17);
  addr_00x_03 <= state_00( 4) & state_00( 0) & state_00(12) & state_00(20);
  addr_00x_04 <= state_00(43) & state_00( 1) & state_00(25) & state_00(19);
  addr_00x_05 <= state_00(16) & state_00(45) & state_00(23) & state_00( 6);
  addr_00x_06 <= state_00(29) & state_00(37) & state_00(11) & state_00(18);
  addr_00x_07 <= state_00(44) & state_00(33) & state_00(42) & state_00(27);
  addr_00x_08 <= state_00( 2) & state_00( 8) & state_00(31) & state_00(47);
  addr_00x_09 <= state_00( 3) & state_00(21) & state_00(28) & state_00( 9);
  addr_00x_10 <= state_00(14) & state_00(35) & state_00(13) & state_00(39);
  addr_00x_11 <= state_00(46) & state_00(30) & state_00( 5) & state_00(22);
  addr_01x_00 <= state_01( 6) & state_01(28) & state_01(16) & state_01(25);
  addr_01x_01 <= state_01( 4) & state_01( 8) & state_01( 0) & state_01(18);
  addr_01x_02 <= state_01(34) & state_01(33) & state_01(37) & state_01(29);
  addr_01x_03 <= state_01(45) & state_01(36) & state_01( 5) & state_01(21);
  addr_01x_04 <= state_01(27) & state_01(13) & state_01(43) & state_01(22);
  addr_01x_05 <= state_01( 2) & state_01(24) & state_01(30) & state_01(42);
  addr_01x_06 <= state_01(12) & state_01(31) & state_01(32) & state_01(10);
  addr_01x_07 <= state_01(46) & state_01(15) & state_01(14) & state_01(47);
  addr_01x_08 <= state_01( 1) & state_01(44) & state_01(19) & state_01(39);
  addr_01x_09 <= state_01( 7) & state_01(38) & state_01(17) & state_01(40);
  addr_01x_10 <= state_01(11) & state_01(26) & state_01(20) & state_01(41);
  addr_01x_11 <= state_01(35) & state_01( 9) & state_01(23) & state_01( 3);
  addr_02x_00 <= state_02(21) & state_02(18) & state_02(12) & state_02(30);
  addr_02x_01 <= state_02(36) & state_02(39) & state_02(44) & state_02(43);
  addr_02x_02 <= state_02(25) & state_02(16) & state_02(35) & state_02(20);
  addr_02x_03 <= state_02( 8) & state_02(11) & state_02( 0) & state_02(15);
  addr_02x_04 <= state_02(14) & state_02(33) & state_02(45) & state_02(41);
  addr_02x_05 <= state_02(27) & state_02( 1) & state_02(38) & state_02(34);
  addr_02x_06 <= state_02(10) & state_02(46) & state_02(47) & state_02(28);
  addr_02x_07 <= state_02( 9) & state_02(29) & state_02(40) & state_02(37);
  addr_02x_08 <= state_02(24) & state_02(19) & state_02( 7) & state_02(22);
  addr_02x_09 <= state_02( 4) & state_02(32) & state_02(13) & state_02(31);
  addr_02x_10 <= state_02( 5) & state_02(42) & state_02( 3) & state_02(23);
  addr_02x_11 <= state_02( 6) & state_02(17) & state_02(26) & state_02( 2);
  addr_03x_00 <= state_03(46) & state_03(47) & state_03(34) & state_03( 9);
  addr_03x_01 <= state_03(37) & state_03(22) & state_03( 2) & state_03(11);
  addr_03x_02 <= state_03( 0) & state_03(39) & state_03(26) & state_03(17);
  addr_03x_03 <= state_03(43) & state_03(10) & state_03(36) & state_03( 7);
  addr_03x_04 <= state_03(32) & state_03(21) & state_03( 3) & state_03( 6);
  addr_03x_05 <= state_03(30) & state_03( 4) & state_03(23) & state_03(40);
  addr_03x_06 <= state_03( 1) & state_03(16) & state_03(38) & state_03(13);
  addr_03x_07 <= state_03(28) & state_03(35) & state_03(19) & state_03(27);
  addr_03x_08 <= state_03(31) & state_03(20) & state_03(12) & state_03(45);
  addr_03x_09 <= state_03(25) & state_03( 8) & state_03(18) & state_03(14);
  addr_03x_10 <= state_03(33) & state_03(44) & state_03(15) & state_03( 5);
  addr_03x_11 <= state_03(24) & state_03(29) & state_03(42) & state_03(41);
  addr_04x_00 <= state_04( 5) & state_04( 7) & state_04(47) & state_04(36);
  addr_04x_01 <= state_04(27) & state_04( 0) & state_04( 6) & state_04(29);
  addr_04x_02 <= state_04(11) & state_04(46) & state_04(39) & state_04(32);
  addr_04x_03 <= state_04(25) & state_04(20) & state_04(10) & state_04(16);
  addr_04x_04 <= state_04(37) & state_04(28) & state_04(30) & state_04(45);
  addr_04x_05 <= state_04( 9) & state_04(22) & state_04(12) & state_04( 1);
  addr_04x_06 <= state_04(38) & state_04(14) & state_04(26) & state_04(18);
  addr_04x_07 <= state_04(44) & state_04(41) & state_04(31) & state_04(24);
  addr_04x_08 <= state_04(35) & state_04(40) & state_04(43) & state_04(17);
  addr_04x_09 <= state_04(33) & state_04(42) & state_04(34) & state_04(13);
  addr_04x_10 <= state_04(21) & state_04(19) & state_04( 2) & state_04(15);
  addr_04x_11 <= state_04(23) & state_04( 4) & state_04( 8) & state_04( 3);
  addr_05x_00 <= state_05(33) & state_05(11) & state_05(30) & state_05( 7);
  addr_05x_01 <= state_05( 5) & state_05(14) & state_05(13) & state_05(27);
  addr_05x_02 <= state_05(47) & state_05(23) & state_05(16) & state_05(39);
  addr_05x_03 <= state_05(31) & state_05(29) & state_05(12) & state_05(41);
  addr_05x_04 <= state_05( 8) & state_05( 1) & state_05(45) & state_05(42);
  addr_05x_05 <= state_05(10) & state_05(36) & state_05( 9) & state_05(15);
  addr_05x_06 <= state_05(32) & state_05(38) & state_05(19) & state_05(40);
  addr_05x_07 <= state_05(43) & state_05(18) & state_05(20) & state_05(34);
  addr_05x_08 <= state_05(26) & state_05( 6) & state_05(46) & state_05( 3);
  addr_05x_09 <= state_05(37) & state_05( 2) & state_05( 4) & state_05(25);
  addr_05x_10 <= state_05(35) & state_05(17) & state_05( 0) & state_05(22);
  addr_05x_11 <= state_05(44) & state_05(28) & state_05(21) & state_05(24);
  addr_06x_00 <= state_06(33) & state_06(10) & state_06(25) & state_06(44);
  addr_06x_01 <= state_06(40) & state_06(24) & state_06(28) & state_06( 2);
  addr_06x_02 <= state_06( 9) & state_06(27) & state_06(17) & state_06( 5);
  addr_06x_03 <= state_06(26) & state_06(14) & state_06( 4) & state_06(22);
  addr_06x_04 <= state_06( 8) & state_06(13) & state_06( 1) & state_06( 3);
  addr_06x_05 <= state_06(41) & state_06(29) & state_06(35) & state_06(42);
  addr_06x_06 <= state_06(34) & state_06(45) & state_06(15) & state_06(20);
  addr_06x_07 <= state_06(18) & state_06(36) & state_06(31) & state_06(32);
  addr_06x_08 <= state_06(39) & state_06(11) & state_06(23) & state_06(19);
  addr_06x_09 <= state_06( 7) & state_06(16) & state_06( 6) & state_06( 0);
  addr_06x_10 <= state_06(21) & state_06(37) & state_06(30) & state_06(46);
  addr_06x_11 <= state_06(43) & state_06(38) & state_06(47) & state_06(12);
  addr_07x_00 <= state_07(22) & state_07(21) & state_07( 9) & state_07(12);
  addr_07x_01 <= state_07(26) & state_07(18) & state_07(41) & state_07(10);
  addr_07x_02 <= state_07(14) & state_07(33) & state_07(39) & state_07(38);
  addr_07x_03 <= state_07(15) & state_07( 3) & state_07(32) & state_07( 6);
  addr_07x_04 <= state_07( 8) & state_07(16) & state_07(31) & state_07(44);
  addr_07x_05 <= state_07(20) & state_07(45) & state_07(40) & state_07(30);
  addr_07x_06 <= state_07( 5) & state_07(34) & state_07(27) & state_07(11);
  addr_07x_07 <= state_07( 7) & state_07(24) & state_07(46) & state_07(13);
  addr_07x_08 <= state_07( 1) & state_07( 2) & state_07(35) & state_07(28);
  addr_07x_09 <= state_07(42) & state_07(17) & state_07(36) & state_07(37);
  addr_07x_10 <= state_07(19) & state_07(23) & state_07(43) & state_07( 0);
  addr_07x_11 <= state_07( 4) & state_07(47) & state_07(25) & state_07(29);
  addr_08x_00 <= state_08(28) & state_08(37) & state_08(33) & state_08( 0);
  addr_08x_01 <= state_08(39) & state_08( 6) & state_08(23) & state_08(41);
  addr_08x_02 <= state_08(35) & state_08(32) & state_08( 3) & state_08(20);
  addr_08x_03 <= state_08(38) & state_08(16) & state_08(17) & state_08(15);
  addr_08x_04 <= state_08(45) & state_08(43) & state_08(36) & state_08(31);
  addr_08x_05 <= state_08(34) & state_08(40) & state_08( 4) & state_08(12);
  addr_08x_06 <= state_08(11) & state_08(47) & state_08(25) & state_08(42);
  addr_08x_07 <= state_08(24) & state_08(14) & state_08( 1) & state_08( 5);
  addr_08x_08 <= state_08(44) & state_08(10) & state_08(27) & state_08( 2);
  addr_08x_09 <= state_08( 9) & state_08(26) & state_08( 8) & state_08(13);
  addr_08x_10 <= state_08(21) & state_08(29) & state_08(46) & state_08(18);
  addr_08x_11 <= state_08(22) & state_08(30) & state_08( 7) & state_08(19);
  addr_09x_00 <= state_09(24) & state_09(17) & state_09(19) & state_09(42);
  addr_09x_01 <= state_09( 9) & state_09(28) & state_09(22) & state_09(25);
  addr_09x_02 <= state_09( 0) & state_09(31) & state_09(46) & state_09(37);
  addr_09x_03 <= state_09(10) & state_09(40) & state_09( 7) & state_09(45);
  addr_09x_04 <= state_09(29) & state_09(11) & state_09(12) & state_09(15);
  addr_09x_05 <= state_09(41) & state_09(13) & state_09( 8) & state_09(36);
  addr_09x_06 <= state_09( 2) & state_09(47) & state_09(35) & state_09( 5);
  addr_09x_07 <= state_09(34) & state_09(18) & state_09(30) & state_09( 1);
  addr_09x_08 <= state_09(27) & state_09(16) & state_09(23) & state_09(43);
  addr_09x_09 <= state_09(32) & state_09( 4) & state_09( 3) & state_09(20);
  addr_09x_10 <= state_09(14) & state_09( 6) & state_09(26) & state_09(38);
  addr_09x_11 <= state_09(44) & state_09(33) & state_09(39) & state_09(21);
  --
  -- State update
  --
  process(enable,clock) is
  begin
    if enable = '1' and rising_edge(clock) then
      -- state 0 update (counter)
      if state_00(23 downto 0) = "101111001101011000001011" then
        carry <= '1';
      else
        carry <= '0';
      end if;
      state_00(23 downto 0) <= std_logic_vector(unsigned(state_00(23 downto 0))+1);
      if carry = '1' then
        state_00(47 downto 24) <= std_logic_vector(unsigned(state_00(47 downto 24))+1);
      end if;
      -- state 1 update (scramble bits using 4x4 S-boxes)
      state_01( 0) <= S_BOX_01_00(to_integer(unsigned(addr_00x_00)));
      state_01( 1) <= S_BOX_01_01(to_integer(unsigned(addr_00x_00)));
      state_01( 2) <= S_BOX_01_02(to_integer(unsigned(addr_00x_00)));
      state_01( 3) <= S_BOX_01_03(to_integer(unsigned(addr_00x_00)));
      state_01( 4) <= S_BOX_01_04(to_integer(unsigned(addr_00x_01)));
      state_01( 5) <= S_BOX_01_05(to_integer(unsigned(addr_00x_01)));
      state_01( 6) <= S_BOX_01_06(to_integer(unsigned(addr_00x_01)));
      state_01( 7) <= S_BOX_01_07(to_integer(unsigned(addr_00x_01)));
      state_01( 8) <= S_BOX_01_08(to_integer(unsigned(addr_00x_02)));
      state_01( 9) <= S_BOX_01_09(to_integer(unsigned(addr_00x_02)));
      state_01(10) <= S_BOX_01_10(to_integer(unsigned(addr_00x_02)));
      state_01(11) <= S_BOX_01_11(to_integer(unsigned(addr_00x_02)));
      state_01(12) <= S_BOX_01_12(to_integer(unsigned(addr_00x_03)));
      state_01(13) <= S_BOX_01_13(to_integer(unsigned(addr_00x_03)));
      state_01(14) <= S_BOX_01_14(to_integer(unsigned(addr_00x_03)));
      state_01(15) <= S_BOX_01_15(to_integer(unsigned(addr_00x_03)));
      state_01(16) <= S_BOX_01_16(to_integer(unsigned(addr_00x_04)));
      state_01(17) <= S_BOX_01_17(to_integer(unsigned(addr_00x_04)));
      state_01(18) <= S_BOX_01_18(to_integer(unsigned(addr_00x_04)));
      state_01(19) <= S_BOX_01_19(to_integer(unsigned(addr_00x_04)));
      state_01(20) <= S_BOX_01_20(to_integer(unsigned(addr_00x_05)));
      state_01(21) <= S_BOX_01_21(to_integer(unsigned(addr_00x_05)));
      state_01(22) <= S_BOX_01_22(to_integer(unsigned(addr_00x_05)));
      state_01(23) <= S_BOX_01_23(to_integer(unsigned(addr_00x_05)));
      state_01(24) <= S_BOX_01_24(to_integer(unsigned(addr_00x_06)));
      state_01(25) <= S_BOX_01_25(to_integer(unsigned(addr_00x_06)));
      state_01(26) <= S_BOX_01_26(to_integer(unsigned(addr_00x_06)));
      state_01(27) <= S_BOX_01_27(to_integer(unsigned(addr_00x_06)));
      state_01(28) <= S_BOX_01_28(to_integer(unsigned(addr_00x_07)));
      state_01(29) <= S_BOX_01_29(to_integer(unsigned(addr_00x_07)));
      state_01(30) <= S_BOX_01_30(to_integer(unsigned(addr_00x_07)));
      state_01(31) <= S_BOX_01_31(to_integer(unsigned(addr_00x_07)));
      state_01(32) <= S_BOX_01_32(to_integer(unsigned(addr_00x_08)));
      state_01(33) <= S_BOX_01_33(to_integer(unsigned(addr_00x_08)));
      state_01(34) <= S_BOX_01_34(to_integer(unsigned(addr_00x_08)));
      state_01(35) <= S_BOX_01_35(to_integer(unsigned(addr_00x_08)));
      state_01(36) <= S_BOX_01_36(to_integer(unsigned(addr_00x_09)));
      state_01(37) <= S_BOX_01_37(to_integer(unsigned(addr_00x_09)));
      state_01(38) <= S_BOX_01_38(to_integer(unsigned(addr_00x_09)));
      state_01(39) <= S_BOX_01_39(to_integer(unsigned(addr_00x_09)));
      state_01(40) <= S_BOX_01_40(to_integer(unsigned(addr_00x_10)));
      state_01(41) <= S_BOX_01_41(to_integer(unsigned(addr_00x_10)));
      state_01(42) <= S_BOX_01_42(to_integer(unsigned(addr_00x_10)));
      state_01(43) <= S_BOX_01_43(to_integer(unsigned(addr_00x_10)));
      state_01(44) <= S_BOX_01_44(to_integer(unsigned(addr_00x_11)));
      state_01(45) <= S_BOX_01_45(to_integer(unsigned(addr_00x_11)));
      state_01(46) <= S_BOX_01_46(to_integer(unsigned(addr_00x_11)));
      state_01(47) <= S_BOX_01_47(to_integer(unsigned(addr_00x_11)));
      -- state 2 update (scramble bits using 4x4 S-boxes)
      state_02( 0) <= S_BOX_02_00(to_integer(unsigned(addr_01x_00)));
      state_02( 1) <= S_BOX_02_01(to_integer(unsigned(addr_01x_00)));
      state_02( 2) <= S_BOX_02_02(to_integer(unsigned(addr_01x_00)));
      state_02( 3) <= S_BOX_02_03(to_integer(unsigned(addr_01x_00)));
      state_02( 4) <= S_BOX_02_04(to_integer(unsigned(addr_01x_01)));
      state_02( 5) <= S_BOX_02_05(to_integer(unsigned(addr_01x_01)));
      state_02( 6) <= S_BOX_02_06(to_integer(unsigned(addr_01x_01)));
      state_02( 7) <= S_BOX_02_07(to_integer(unsigned(addr_01x_01)));
      state_02( 8) <= S_BOX_02_08(to_integer(unsigned(addr_01x_02)));
      state_02( 9) <= S_BOX_02_09(to_integer(unsigned(addr_01x_02)));
      state_02(10) <= S_BOX_02_10(to_integer(unsigned(addr_01x_02)));
      state_02(11) <= S_BOX_02_11(to_integer(unsigned(addr_01x_02)));
      state_02(12) <= S_BOX_02_12(to_integer(unsigned(addr_01x_03)));
      state_02(13) <= S_BOX_02_13(to_integer(unsigned(addr_01x_03)));
      state_02(14) <= S_BOX_02_14(to_integer(unsigned(addr_01x_03)));
      state_02(15) <= S_BOX_02_15(to_integer(unsigned(addr_01x_03)));
      state_02(16) <= S_BOX_02_16(to_integer(unsigned(addr_01x_04)));
      state_02(17) <= S_BOX_02_17(to_integer(unsigned(addr_01x_04)));
      state_02(18) <= S_BOX_02_18(to_integer(unsigned(addr_01x_04)));
      state_02(19) <= S_BOX_02_19(to_integer(unsigned(addr_01x_04)));
      state_02(20) <= S_BOX_02_20(to_integer(unsigned(addr_01x_05)));
      state_02(21) <= S_BOX_02_21(to_integer(unsigned(addr_01x_05)));
      state_02(22) <= S_BOX_02_22(to_integer(unsigned(addr_01x_05)));
      state_02(23) <= S_BOX_02_23(to_integer(unsigned(addr_01x_05)));
      state_02(24) <= S_BOX_02_24(to_integer(unsigned(addr_01x_06)));
      state_02(25) <= S_BOX_02_25(to_integer(unsigned(addr_01x_06)));
      state_02(26) <= S_BOX_02_26(to_integer(unsigned(addr_01x_06)));
      state_02(27) <= S_BOX_02_27(to_integer(unsigned(addr_01x_06)));
      state_02(28) <= S_BOX_02_28(to_integer(unsigned(addr_01x_07)));
      state_02(29) <= S_BOX_02_29(to_integer(unsigned(addr_01x_07)));
      state_02(30) <= S_BOX_02_30(to_integer(unsigned(addr_01x_07)));
      state_02(31) <= S_BOX_02_31(to_integer(unsigned(addr_01x_07)));
      state_02(32) <= S_BOX_02_32(to_integer(unsigned(addr_01x_08)));
      state_02(33) <= S_BOX_02_33(to_integer(unsigned(addr_01x_08)));
      state_02(34) <= S_BOX_02_34(to_integer(unsigned(addr_01x_08)));
      state_02(35) <= S_BOX_02_35(to_integer(unsigned(addr_01x_08)));
      state_02(36) <= S_BOX_02_36(to_integer(unsigned(addr_01x_09)));
      state_02(37) <= S_BOX_02_37(to_integer(unsigned(addr_01x_09)));
      state_02(38) <= S_BOX_02_38(to_integer(unsigned(addr_01x_09)));
      state_02(39) <= S_BOX_02_39(to_integer(unsigned(addr_01x_09)));
      state_02(40) <= S_BOX_02_40(to_integer(unsigned(addr_01x_10)));
      state_02(41) <= S_BOX_02_41(to_integer(unsigned(addr_01x_10)));
      state_02(42) <= S_BOX_02_42(to_integer(unsigned(addr_01x_10)));
      state_02(43) <= S_BOX_02_43(to_integer(unsigned(addr_01x_10)));
      state_02(44) <= S_BOX_02_44(to_integer(unsigned(addr_01x_11)));
      state_02(45) <= S_BOX_02_45(to_integer(unsigned(addr_01x_11)));
      state_02(46) <= S_BOX_02_46(to_integer(unsigned(addr_01x_11)));
      state_02(47) <= S_BOX_02_47(to_integer(unsigned(addr_01x_11)));
      -- state 3 update (scramble bits using 4x4 S-boxes)
      state_03( 0) <= S_BOX_03_00(to_integer(unsigned(addr_02x_00)));
      state_03( 1) <= S_BOX_03_01(to_integer(unsigned(addr_02x_00)));
      state_03( 2) <= S_BOX_03_02(to_integer(unsigned(addr_02x_00)));
      state_03( 3) <= S_BOX_03_03(to_integer(unsigned(addr_02x_00)));
      state_03( 4) <= S_BOX_03_04(to_integer(unsigned(addr_02x_01)));
      state_03( 5) <= S_BOX_03_05(to_integer(unsigned(addr_02x_01)));
      state_03( 6) <= S_BOX_03_06(to_integer(unsigned(addr_02x_01)));
      state_03( 7) <= S_BOX_03_07(to_integer(unsigned(addr_02x_01)));
      state_03( 8) <= S_BOX_03_08(to_integer(unsigned(addr_02x_02)));
      state_03( 9) <= S_BOX_03_09(to_integer(unsigned(addr_02x_02)));
      state_03(10) <= S_BOX_03_10(to_integer(unsigned(addr_02x_02)));
      state_03(11) <= S_BOX_03_11(to_integer(unsigned(addr_02x_02)));
      state_03(12) <= S_BOX_03_12(to_integer(unsigned(addr_02x_03)));
      state_03(13) <= S_BOX_03_13(to_integer(unsigned(addr_02x_03)));
      state_03(14) <= S_BOX_03_14(to_integer(unsigned(addr_02x_03)));
      state_03(15) <= S_BOX_03_15(to_integer(unsigned(addr_02x_03)));
      state_03(16) <= S_BOX_03_16(to_integer(unsigned(addr_02x_04)));
      state_03(17) <= S_BOX_03_17(to_integer(unsigned(addr_02x_04)));
      state_03(18) <= S_BOX_03_18(to_integer(unsigned(addr_02x_04)));
      state_03(19) <= S_BOX_03_19(to_integer(unsigned(addr_02x_04)));
      state_03(20) <= S_BOX_03_20(to_integer(unsigned(addr_02x_05)));
      state_03(21) <= S_BOX_03_21(to_integer(unsigned(addr_02x_05)));
      state_03(22) <= S_BOX_03_22(to_integer(unsigned(addr_02x_05)));
      state_03(23) <= S_BOX_03_23(to_integer(unsigned(addr_02x_05)));
      state_03(24) <= S_BOX_03_24(to_integer(unsigned(addr_02x_06)));
      state_03(25) <= S_BOX_03_25(to_integer(unsigned(addr_02x_06)));
      state_03(26) <= S_BOX_03_26(to_integer(unsigned(addr_02x_06)));
      state_03(27) <= S_BOX_03_27(to_integer(unsigned(addr_02x_06)));
      state_03(28) <= S_BOX_03_28(to_integer(unsigned(addr_02x_07)));
      state_03(29) <= S_BOX_03_29(to_integer(unsigned(addr_02x_07)));
      state_03(30) <= S_BOX_03_30(to_integer(unsigned(addr_02x_07)));
      state_03(31) <= S_BOX_03_31(to_integer(unsigned(addr_02x_07)));
      state_03(32) <= S_BOX_03_32(to_integer(unsigned(addr_02x_08)));
      state_03(33) <= S_BOX_03_33(to_integer(unsigned(addr_02x_08)));
      state_03(34) <= S_BOX_03_34(to_integer(unsigned(addr_02x_08)));
      state_03(35) <= S_BOX_03_35(to_integer(unsigned(addr_02x_08)));
      state_03(36) <= S_BOX_03_36(to_integer(unsigned(addr_02x_09)));
      state_03(37) <= S_BOX_03_37(to_integer(unsigned(addr_02x_09)));
      state_03(38) <= S_BOX_03_38(to_integer(unsigned(addr_02x_09)));
      state_03(39) <= S_BOX_03_39(to_integer(unsigned(addr_02x_09)));
      state_03(40) <= S_BOX_03_40(to_integer(unsigned(addr_02x_10)));
      state_03(41) <= S_BOX_03_41(to_integer(unsigned(addr_02x_10)));
      state_03(42) <= S_BOX_03_42(to_integer(unsigned(addr_02x_10)));
      state_03(43) <= S_BOX_03_43(to_integer(unsigned(addr_02x_10)));
      state_03(44) <= S_BOX_03_44(to_integer(unsigned(addr_02x_11)));
      state_03(45) <= S_BOX_03_45(to_integer(unsigned(addr_02x_11)));
      state_03(46) <= S_BOX_03_46(to_integer(unsigned(addr_02x_11)));
      state_03(47) <= S_BOX_03_47(to_integer(unsigned(addr_02x_11)));
      -- state 4 update (scramble bits using 4x4 S-boxes)
      state_04( 0) <= S_BOX_04_00(to_integer(unsigned(addr_03x_00)));
      state_04( 1) <= S_BOX_04_01(to_integer(unsigned(addr_03x_00)));
      state_04( 2) <= S_BOX_04_02(to_integer(unsigned(addr_03x_00)));
      state_04( 3) <= S_BOX_04_03(to_integer(unsigned(addr_03x_00)));
      state_04( 4) <= S_BOX_04_04(to_integer(unsigned(addr_03x_01)));
      state_04( 5) <= S_BOX_04_05(to_integer(unsigned(addr_03x_01)));
      state_04( 6) <= S_BOX_04_06(to_integer(unsigned(addr_03x_01)));
      state_04( 7) <= S_BOX_04_07(to_integer(unsigned(addr_03x_01)));
      state_04( 8) <= S_BOX_04_08(to_integer(unsigned(addr_03x_02)));
      state_04( 9) <= S_BOX_04_09(to_integer(unsigned(addr_03x_02)));
      state_04(10) <= S_BOX_04_10(to_integer(unsigned(addr_03x_02)));
      state_04(11) <= S_BOX_04_11(to_integer(unsigned(addr_03x_02)));
      state_04(12) <= S_BOX_04_12(to_integer(unsigned(addr_03x_03)));
      state_04(13) <= S_BOX_04_13(to_integer(unsigned(addr_03x_03)));
      state_04(14) <= S_BOX_04_14(to_integer(unsigned(addr_03x_03)));
      state_04(15) <= S_BOX_04_15(to_integer(unsigned(addr_03x_03)));
      state_04(16) <= S_BOX_04_16(to_integer(unsigned(addr_03x_04)));
      state_04(17) <= S_BOX_04_17(to_integer(unsigned(addr_03x_04)));
      state_04(18) <= S_BOX_04_18(to_integer(unsigned(addr_03x_04)));
      state_04(19) <= S_BOX_04_19(to_integer(unsigned(addr_03x_04)));
      state_04(20) <= S_BOX_04_20(to_integer(unsigned(addr_03x_05)));
      state_04(21) <= S_BOX_04_21(to_integer(unsigned(addr_03x_05)));
      state_04(22) <= S_BOX_04_22(to_integer(unsigned(addr_03x_05)));
      state_04(23) <= S_BOX_04_23(to_integer(unsigned(addr_03x_05)));
      state_04(24) <= S_BOX_04_24(to_integer(unsigned(addr_03x_06)));
      state_04(25) <= S_BOX_04_25(to_integer(unsigned(addr_03x_06)));
      state_04(26) <= S_BOX_04_26(to_integer(unsigned(addr_03x_06)));
      state_04(27) <= S_BOX_04_27(to_integer(unsigned(addr_03x_06)));
      state_04(28) <= S_BOX_04_28(to_integer(unsigned(addr_03x_07)));
      state_04(29) <= S_BOX_04_29(to_integer(unsigned(addr_03x_07)));
      state_04(30) <= S_BOX_04_30(to_integer(unsigned(addr_03x_07)));
      state_04(31) <= S_BOX_04_31(to_integer(unsigned(addr_03x_07)));
      state_04(32) <= S_BOX_04_32(to_integer(unsigned(addr_03x_08)));
      state_04(33) <= S_BOX_04_33(to_integer(unsigned(addr_03x_08)));
      state_04(34) <= S_BOX_04_34(to_integer(unsigned(addr_03x_08)));
      state_04(35) <= S_BOX_04_35(to_integer(unsigned(addr_03x_08)));
      state_04(36) <= S_BOX_04_36(to_integer(unsigned(addr_03x_09)));
      state_04(37) <= S_BOX_04_37(to_integer(unsigned(addr_03x_09)));
      state_04(38) <= S_BOX_04_38(to_integer(unsigned(addr_03x_09)));
      state_04(39) <= S_BOX_04_39(to_integer(unsigned(addr_03x_09)));
      state_04(40) <= S_BOX_04_40(to_integer(unsigned(addr_03x_10)));
      state_04(41) <= S_BOX_04_41(to_integer(unsigned(addr_03x_10)));
      state_04(42) <= S_BOX_04_42(to_integer(unsigned(addr_03x_10)));
      state_04(43) <= S_BOX_04_43(to_integer(unsigned(addr_03x_10)));
      state_04(44) <= S_BOX_04_44(to_integer(unsigned(addr_03x_11)));
      state_04(45) <= S_BOX_04_45(to_integer(unsigned(addr_03x_11)));
      state_04(46) <= S_BOX_04_46(to_integer(unsigned(addr_03x_11)));
      state_04(47) <= S_BOX_04_47(to_integer(unsigned(addr_03x_11)));
      -- state 5 update (scramble bits using 4x4 S-boxes)
      state_05( 0) <= S_BOX_05_00(to_integer(unsigned(addr_04x_00)));
      state_05( 1) <= S_BOX_05_01(to_integer(unsigned(addr_04x_00)));
      state_05( 2) <= S_BOX_05_02(to_integer(unsigned(addr_04x_00)));
      state_05( 3) <= S_BOX_05_03(to_integer(unsigned(addr_04x_00)));
      state_05( 4) <= S_BOX_05_04(to_integer(unsigned(addr_04x_01)));
      state_05( 5) <= S_BOX_05_05(to_integer(unsigned(addr_04x_01)));
      state_05( 6) <= S_BOX_05_06(to_integer(unsigned(addr_04x_01)));
      state_05( 7) <= S_BOX_05_07(to_integer(unsigned(addr_04x_01)));
      state_05( 8) <= S_BOX_05_08(to_integer(unsigned(addr_04x_02)));
      state_05( 9) <= S_BOX_05_09(to_integer(unsigned(addr_04x_02)));
      state_05(10) <= S_BOX_05_10(to_integer(unsigned(addr_04x_02)));
      state_05(11) <= S_BOX_05_11(to_integer(unsigned(addr_04x_02)));
      state_05(12) <= S_BOX_05_12(to_integer(unsigned(addr_04x_03)));
      state_05(13) <= S_BOX_05_13(to_integer(unsigned(addr_04x_03)));
      state_05(14) <= S_BOX_05_14(to_integer(unsigned(addr_04x_03)));
      state_05(15) <= S_BOX_05_15(to_integer(unsigned(addr_04x_03)));
      state_05(16) <= S_BOX_05_16(to_integer(unsigned(addr_04x_04)));
      state_05(17) <= S_BOX_05_17(to_integer(unsigned(addr_04x_04)));
      state_05(18) <= S_BOX_05_18(to_integer(unsigned(addr_04x_04)));
      state_05(19) <= S_BOX_05_19(to_integer(unsigned(addr_04x_04)));
      state_05(20) <= S_BOX_05_20(to_integer(unsigned(addr_04x_05)));
      state_05(21) <= S_BOX_05_21(to_integer(unsigned(addr_04x_05)));
      state_05(22) <= S_BOX_05_22(to_integer(unsigned(addr_04x_05)));
      state_05(23) <= S_BOX_05_23(to_integer(unsigned(addr_04x_05)));
      state_05(24) <= S_BOX_05_24(to_integer(unsigned(addr_04x_06)));
      state_05(25) <= S_BOX_05_25(to_integer(unsigned(addr_04x_06)));
      state_05(26) <= S_BOX_05_26(to_integer(unsigned(addr_04x_06)));
      state_05(27) <= S_BOX_05_27(to_integer(unsigned(addr_04x_06)));
      state_05(28) <= S_BOX_05_28(to_integer(unsigned(addr_04x_07)));
      state_05(29) <= S_BOX_05_29(to_integer(unsigned(addr_04x_07)));
      state_05(30) <= S_BOX_05_30(to_integer(unsigned(addr_04x_07)));
      state_05(31) <= S_BOX_05_31(to_integer(unsigned(addr_04x_07)));
      state_05(32) <= S_BOX_05_32(to_integer(unsigned(addr_04x_08)));
      state_05(33) <= S_BOX_05_33(to_integer(unsigned(addr_04x_08)));
      state_05(34) <= S_BOX_05_34(to_integer(unsigned(addr_04x_08)));
      state_05(35) <= S_BOX_05_35(to_integer(unsigned(addr_04x_08)));
      state_05(36) <= S_BOX_05_36(to_integer(unsigned(addr_04x_09)));
      state_05(37) <= S_BOX_05_37(to_integer(unsigned(addr_04x_09)));
      state_05(38) <= S_BOX_05_38(to_integer(unsigned(addr_04x_09)));
      state_05(39) <= S_BOX_05_39(to_integer(unsigned(addr_04x_09)));
      state_05(40) <= S_BOX_05_40(to_integer(unsigned(addr_04x_10)));
      state_05(41) <= S_BOX_05_41(to_integer(unsigned(addr_04x_10)));
      state_05(42) <= S_BOX_05_42(to_integer(unsigned(addr_04x_10)));
      state_05(43) <= S_BOX_05_43(to_integer(unsigned(addr_04x_10)));
      state_05(44) <= S_BOX_05_44(to_integer(unsigned(addr_04x_11)));
      state_05(45) <= S_BOX_05_45(to_integer(unsigned(addr_04x_11)));
      state_05(46) <= S_BOX_05_46(to_integer(unsigned(addr_04x_11)));
      state_05(47) <= S_BOX_05_47(to_integer(unsigned(addr_04x_11)));
      -- state 6 update (scramble bits using 4x4 S-boxes)
      state_06( 0) <= S_BOX_06_00(to_integer(unsigned(addr_05x_00)));
      state_06( 1) <= S_BOX_06_01(to_integer(unsigned(addr_05x_00)));
      state_06( 2) <= S_BOX_06_02(to_integer(unsigned(addr_05x_00)));
      state_06( 3) <= S_BOX_06_03(to_integer(unsigned(addr_05x_00)));
      state_06( 4) <= S_BOX_06_04(to_integer(unsigned(addr_05x_01)));
      state_06( 5) <= S_BOX_06_05(to_integer(unsigned(addr_05x_01)));
      state_06( 6) <= S_BOX_06_06(to_integer(unsigned(addr_05x_01)));
      state_06( 7) <= S_BOX_06_07(to_integer(unsigned(addr_05x_01)));
      state_06( 8) <= S_BOX_06_08(to_integer(unsigned(addr_05x_02)));
      state_06( 9) <= S_BOX_06_09(to_integer(unsigned(addr_05x_02)));
      state_06(10) <= S_BOX_06_10(to_integer(unsigned(addr_05x_02)));
      state_06(11) <= S_BOX_06_11(to_integer(unsigned(addr_05x_02)));
      state_06(12) <= S_BOX_06_12(to_integer(unsigned(addr_05x_03)));
      state_06(13) <= S_BOX_06_13(to_integer(unsigned(addr_05x_03)));
      state_06(14) <= S_BOX_06_14(to_integer(unsigned(addr_05x_03)));
      state_06(15) <= S_BOX_06_15(to_integer(unsigned(addr_05x_03)));
      state_06(16) <= S_BOX_06_16(to_integer(unsigned(addr_05x_04)));
      state_06(17) <= S_BOX_06_17(to_integer(unsigned(addr_05x_04)));
      state_06(18) <= S_BOX_06_18(to_integer(unsigned(addr_05x_04)));
      state_06(19) <= S_BOX_06_19(to_integer(unsigned(addr_05x_04)));
      state_06(20) <= S_BOX_06_20(to_integer(unsigned(addr_05x_05)));
      state_06(21) <= S_BOX_06_21(to_integer(unsigned(addr_05x_05)));
      state_06(22) <= S_BOX_06_22(to_integer(unsigned(addr_05x_05)));
      state_06(23) <= S_BOX_06_23(to_integer(unsigned(addr_05x_05)));
      state_06(24) <= S_BOX_06_24(to_integer(unsigned(addr_05x_06)));
      state_06(25) <= S_BOX_06_25(to_integer(unsigned(addr_05x_06)));
      state_06(26) <= S_BOX_06_26(to_integer(unsigned(addr_05x_06)));
      state_06(27) <= S_BOX_06_27(to_integer(unsigned(addr_05x_06)));
      state_06(28) <= S_BOX_06_28(to_integer(unsigned(addr_05x_07)));
      state_06(29) <= S_BOX_06_29(to_integer(unsigned(addr_05x_07)));
      state_06(30) <= S_BOX_06_30(to_integer(unsigned(addr_05x_07)));
      state_06(31) <= S_BOX_06_31(to_integer(unsigned(addr_05x_07)));
      state_06(32) <= S_BOX_06_32(to_integer(unsigned(addr_05x_08)));
      state_06(33) <= S_BOX_06_33(to_integer(unsigned(addr_05x_08)));
      state_06(34) <= S_BOX_06_34(to_integer(unsigned(addr_05x_08)));
      state_06(35) <= S_BOX_06_35(to_integer(unsigned(addr_05x_08)));
      state_06(36) <= S_BOX_06_36(to_integer(unsigned(addr_05x_09)));
      state_06(37) <= S_BOX_06_37(to_integer(unsigned(addr_05x_09)));
      state_06(38) <= S_BOX_06_38(to_integer(unsigned(addr_05x_09)));
      state_06(39) <= S_BOX_06_39(to_integer(unsigned(addr_05x_09)));
      state_06(40) <= S_BOX_06_40(to_integer(unsigned(addr_05x_10)));
      state_06(41) <= S_BOX_06_41(to_integer(unsigned(addr_05x_10)));
      state_06(42) <= S_BOX_06_42(to_integer(unsigned(addr_05x_10)));
      state_06(43) <= S_BOX_06_43(to_integer(unsigned(addr_05x_10)));
      state_06(44) <= S_BOX_06_44(to_integer(unsigned(addr_05x_11)));
      state_06(45) <= S_BOX_06_45(to_integer(unsigned(addr_05x_11)));
      state_06(46) <= S_BOX_06_46(to_integer(unsigned(addr_05x_11)));
      state_06(47) <= S_BOX_06_47(to_integer(unsigned(addr_05x_11)));
      -- state 7 update (scramble bits using 4x4 S-boxes)
      state_07( 0) <= S_BOX_07_00(to_integer(unsigned(addr_06x_00)));
      state_07( 1) <= S_BOX_07_01(to_integer(unsigned(addr_06x_00)));
      state_07( 2) <= S_BOX_07_02(to_integer(unsigned(addr_06x_00)));
      state_07( 3) <= S_BOX_07_03(to_integer(unsigned(addr_06x_00)));
      state_07( 4) <= S_BOX_07_04(to_integer(unsigned(addr_06x_01)));
      state_07( 5) <= S_BOX_07_05(to_integer(unsigned(addr_06x_01)));
      state_07( 6) <= S_BOX_07_06(to_integer(unsigned(addr_06x_01)));
      state_07( 7) <= S_BOX_07_07(to_integer(unsigned(addr_06x_01)));
      state_07( 8) <= S_BOX_07_08(to_integer(unsigned(addr_06x_02)));
      state_07( 9) <= S_BOX_07_09(to_integer(unsigned(addr_06x_02)));
      state_07(10) <= S_BOX_07_10(to_integer(unsigned(addr_06x_02)));
      state_07(11) <= S_BOX_07_11(to_integer(unsigned(addr_06x_02)));
      state_07(12) <= S_BOX_07_12(to_integer(unsigned(addr_06x_03)));
      state_07(13) <= S_BOX_07_13(to_integer(unsigned(addr_06x_03)));
      state_07(14) <= S_BOX_07_14(to_integer(unsigned(addr_06x_03)));
      state_07(15) <= S_BOX_07_15(to_integer(unsigned(addr_06x_03)));
      state_07(16) <= S_BOX_07_16(to_integer(unsigned(addr_06x_04)));
      state_07(17) <= S_BOX_07_17(to_integer(unsigned(addr_06x_04)));
      state_07(18) <= S_BOX_07_18(to_integer(unsigned(addr_06x_04)));
      state_07(19) <= S_BOX_07_19(to_integer(unsigned(addr_06x_04)));
      state_07(20) <= S_BOX_07_20(to_integer(unsigned(addr_06x_05)));
      state_07(21) <= S_BOX_07_21(to_integer(unsigned(addr_06x_05)));
      state_07(22) <= S_BOX_07_22(to_integer(unsigned(addr_06x_05)));
      state_07(23) <= S_BOX_07_23(to_integer(unsigned(addr_06x_05)));
      state_07(24) <= S_BOX_07_24(to_integer(unsigned(addr_06x_06)));
      state_07(25) <= S_BOX_07_25(to_integer(unsigned(addr_06x_06)));
      state_07(26) <= S_BOX_07_26(to_integer(unsigned(addr_06x_06)));
      state_07(27) <= S_BOX_07_27(to_integer(unsigned(addr_06x_06)));
      state_07(28) <= S_BOX_07_28(to_integer(unsigned(addr_06x_07)));
      state_07(29) <= S_BOX_07_29(to_integer(unsigned(addr_06x_07)));
      state_07(30) <= S_BOX_07_30(to_integer(unsigned(addr_06x_07)));
      state_07(31) <= S_BOX_07_31(to_integer(unsigned(addr_06x_07)));
      state_07(32) <= S_BOX_07_32(to_integer(unsigned(addr_06x_08)));
      state_07(33) <= S_BOX_07_33(to_integer(unsigned(addr_06x_08)));
      state_07(34) <= S_BOX_07_34(to_integer(unsigned(addr_06x_08)));
      state_07(35) <= S_BOX_07_35(to_integer(unsigned(addr_06x_08)));
      state_07(36) <= S_BOX_07_36(to_integer(unsigned(addr_06x_09)));
      state_07(37) <= S_BOX_07_37(to_integer(unsigned(addr_06x_09)));
      state_07(38) <= S_BOX_07_38(to_integer(unsigned(addr_06x_09)));
      state_07(39) <= S_BOX_07_39(to_integer(unsigned(addr_06x_09)));
      state_07(40) <= S_BOX_07_40(to_integer(unsigned(addr_06x_10)));
      state_07(41) <= S_BOX_07_41(to_integer(unsigned(addr_06x_10)));
      state_07(42) <= S_BOX_07_42(to_integer(unsigned(addr_06x_10)));
      state_07(43) <= S_BOX_07_43(to_integer(unsigned(addr_06x_10)));
      state_07(44) <= S_BOX_07_44(to_integer(unsigned(addr_06x_11)));
      state_07(45) <= S_BOX_07_45(to_integer(unsigned(addr_06x_11)));
      state_07(46) <= S_BOX_07_46(to_integer(unsigned(addr_06x_11)));
      state_07(47) <= S_BOX_07_47(to_integer(unsigned(addr_06x_11)));
      -- state 8 update (scramble bits using 4x4 S-boxes)
      state_08( 0) <= S_BOX_08_00(to_integer(unsigned(addr_07x_00)));
      state_08( 1) <= S_BOX_08_01(to_integer(unsigned(addr_07x_00)));
      state_08( 2) <= S_BOX_08_02(to_integer(unsigned(addr_07x_00)));
      state_08( 3) <= S_BOX_08_03(to_integer(unsigned(addr_07x_00)));
      state_08( 4) <= S_BOX_08_04(to_integer(unsigned(addr_07x_01)));
      state_08( 5) <= S_BOX_08_05(to_integer(unsigned(addr_07x_01)));
      state_08( 6) <= S_BOX_08_06(to_integer(unsigned(addr_07x_01)));
      state_08( 7) <= S_BOX_08_07(to_integer(unsigned(addr_07x_01)));
      state_08( 8) <= S_BOX_08_08(to_integer(unsigned(addr_07x_02)));
      state_08( 9) <= S_BOX_08_09(to_integer(unsigned(addr_07x_02)));
      state_08(10) <= S_BOX_08_10(to_integer(unsigned(addr_07x_02)));
      state_08(11) <= S_BOX_08_11(to_integer(unsigned(addr_07x_02)));
      state_08(12) <= S_BOX_08_12(to_integer(unsigned(addr_07x_03)));
      state_08(13) <= S_BOX_08_13(to_integer(unsigned(addr_07x_03)));
      state_08(14) <= S_BOX_08_14(to_integer(unsigned(addr_07x_03)));
      state_08(15) <= S_BOX_08_15(to_integer(unsigned(addr_07x_03)));
      state_08(16) <= S_BOX_08_16(to_integer(unsigned(addr_07x_04)));
      state_08(17) <= S_BOX_08_17(to_integer(unsigned(addr_07x_04)));
      state_08(18) <= S_BOX_08_18(to_integer(unsigned(addr_07x_04)));
      state_08(19) <= S_BOX_08_19(to_integer(unsigned(addr_07x_04)));
      state_08(20) <= S_BOX_08_20(to_integer(unsigned(addr_07x_05)));
      state_08(21) <= S_BOX_08_21(to_integer(unsigned(addr_07x_05)));
      state_08(22) <= S_BOX_08_22(to_integer(unsigned(addr_07x_05)));
      state_08(23) <= S_BOX_08_23(to_integer(unsigned(addr_07x_05)));
      state_08(24) <= S_BOX_08_24(to_integer(unsigned(addr_07x_06)));
      state_08(25) <= S_BOX_08_25(to_integer(unsigned(addr_07x_06)));
      state_08(26) <= S_BOX_08_26(to_integer(unsigned(addr_07x_06)));
      state_08(27) <= S_BOX_08_27(to_integer(unsigned(addr_07x_06)));
      state_08(28) <= S_BOX_08_28(to_integer(unsigned(addr_07x_07)));
      state_08(29) <= S_BOX_08_29(to_integer(unsigned(addr_07x_07)));
      state_08(30) <= S_BOX_08_30(to_integer(unsigned(addr_07x_07)));
      state_08(31) <= S_BOX_08_31(to_integer(unsigned(addr_07x_07)));
      state_08(32) <= S_BOX_08_32(to_integer(unsigned(addr_07x_08)));
      state_08(33) <= S_BOX_08_33(to_integer(unsigned(addr_07x_08)));
      state_08(34) <= S_BOX_08_34(to_integer(unsigned(addr_07x_08)));
      state_08(35) <= S_BOX_08_35(to_integer(unsigned(addr_07x_08)));
      state_08(36) <= S_BOX_08_36(to_integer(unsigned(addr_07x_09)));
      state_08(37) <= S_BOX_08_37(to_integer(unsigned(addr_07x_09)));
      state_08(38) <= S_BOX_08_38(to_integer(unsigned(addr_07x_09)));
      state_08(39) <= S_BOX_08_39(to_integer(unsigned(addr_07x_09)));
      state_08(40) <= S_BOX_08_40(to_integer(unsigned(addr_07x_10)));
      state_08(41) <= S_BOX_08_41(to_integer(unsigned(addr_07x_10)));
      state_08(42) <= S_BOX_08_42(to_integer(unsigned(addr_07x_10)));
      state_08(43) <= S_BOX_08_43(to_integer(unsigned(addr_07x_10)));
      state_08(44) <= S_BOX_08_44(to_integer(unsigned(addr_07x_11)));
      state_08(45) <= S_BOX_08_45(to_integer(unsigned(addr_07x_11)));
      state_08(46) <= S_BOX_08_46(to_integer(unsigned(addr_07x_11)));
      state_08(47) <= S_BOX_08_47(to_integer(unsigned(addr_07x_11)));
      -- state 9 update (scramble bits using 4x4 S-boxes)
      state_09( 0) <= S_BOX_09_00(to_integer(unsigned(addr_08x_00)));
      state_09( 1) <= S_BOX_09_01(to_integer(unsigned(addr_08x_00)));
      state_09( 2) <= S_BOX_09_02(to_integer(unsigned(addr_08x_00)));
      state_09( 3) <= S_BOX_09_03(to_integer(unsigned(addr_08x_00)));
      state_09( 4) <= S_BOX_09_04(to_integer(unsigned(addr_08x_01)));
      state_09( 5) <= S_BOX_09_05(to_integer(unsigned(addr_08x_01)));
      state_09( 6) <= S_BOX_09_06(to_integer(unsigned(addr_08x_01)));
      state_09( 7) <= S_BOX_09_07(to_integer(unsigned(addr_08x_01)));
      state_09( 8) <= S_BOX_09_08(to_integer(unsigned(addr_08x_02)));
      state_09( 9) <= S_BOX_09_09(to_integer(unsigned(addr_08x_02)));
      state_09(10) <= S_BOX_09_10(to_integer(unsigned(addr_08x_02)));
      state_09(11) <= S_BOX_09_11(to_integer(unsigned(addr_08x_02)));
      state_09(12) <= S_BOX_09_12(to_integer(unsigned(addr_08x_03)));
      state_09(13) <= S_BOX_09_13(to_integer(unsigned(addr_08x_03)));
      state_09(14) <= S_BOX_09_14(to_integer(unsigned(addr_08x_03)));
      state_09(15) <= S_BOX_09_15(to_integer(unsigned(addr_08x_03)));
      state_09(16) <= S_BOX_09_16(to_integer(unsigned(addr_08x_04)));
      state_09(17) <= S_BOX_09_17(to_integer(unsigned(addr_08x_04)));
      state_09(18) <= S_BOX_09_18(to_integer(unsigned(addr_08x_04)));
      state_09(19) <= S_BOX_09_19(to_integer(unsigned(addr_08x_04)));
      state_09(20) <= S_BOX_09_20(to_integer(unsigned(addr_08x_05)));
      state_09(21) <= S_BOX_09_21(to_integer(unsigned(addr_08x_05)));
      state_09(22) <= S_BOX_09_22(to_integer(unsigned(addr_08x_05)));
      state_09(23) <= S_BOX_09_23(to_integer(unsigned(addr_08x_05)));
      state_09(24) <= S_BOX_09_24(to_integer(unsigned(addr_08x_06)));
      state_09(25) <= S_BOX_09_25(to_integer(unsigned(addr_08x_06)));
      state_09(26) <= S_BOX_09_26(to_integer(unsigned(addr_08x_06)));
      state_09(27) <= S_BOX_09_27(to_integer(unsigned(addr_08x_06)));
      state_09(28) <= S_BOX_09_28(to_integer(unsigned(addr_08x_07)));
      state_09(29) <= S_BOX_09_29(to_integer(unsigned(addr_08x_07)));
      state_09(30) <= S_BOX_09_30(to_integer(unsigned(addr_08x_07)));
      state_09(31) <= S_BOX_09_31(to_integer(unsigned(addr_08x_07)));
      state_09(32) <= S_BOX_09_32(to_integer(unsigned(addr_08x_08)));
      state_09(33) <= S_BOX_09_33(to_integer(unsigned(addr_08x_08)));
      state_09(34) <= S_BOX_09_34(to_integer(unsigned(addr_08x_08)));
      state_09(35) <= S_BOX_09_35(to_integer(unsigned(addr_08x_08)));
      state_09(36) <= S_BOX_09_36(to_integer(unsigned(addr_08x_09)));
      state_09(37) <= S_BOX_09_37(to_integer(unsigned(addr_08x_09)));
      state_09(38) <= S_BOX_09_38(to_integer(unsigned(addr_08x_09)));
      state_09(39) <= S_BOX_09_39(to_integer(unsigned(addr_08x_09)));
      state_09(40) <= S_BOX_09_40(to_integer(unsigned(addr_08x_10)));
      state_09(41) <= S_BOX_09_41(to_integer(unsigned(addr_08x_10)));
      state_09(42) <= S_BOX_09_42(to_integer(unsigned(addr_08x_10)));
      state_09(43) <= S_BOX_09_43(to_integer(unsigned(addr_08x_10)));
      state_09(44) <= S_BOX_09_44(to_integer(unsigned(addr_08x_11)));
      state_09(45) <= S_BOX_09_45(to_integer(unsigned(addr_08x_11)));
      state_09(46) <= S_BOX_09_46(to_integer(unsigned(addr_08x_11)));
      state_09(47) <= S_BOX_09_47(to_integer(unsigned(addr_08x_11)));
      -- state 10 update (scramble bits using 4x4 S-boxes)
      state_10( 0) <= S_BOX_10_00(to_integer(unsigned(addr_09x_00)));
      state_10( 1) <= S_BOX_10_01(to_integer(unsigned(addr_09x_00)));
      state_10( 2) <= S_BOX_10_02(to_integer(unsigned(addr_09x_00)));
      state_10( 3) <= S_BOX_10_03(to_integer(unsigned(addr_09x_00)));
      state_10( 4) <= S_BOX_10_04(to_integer(unsigned(addr_09x_01)));
      state_10( 5) <= S_BOX_10_05(to_integer(unsigned(addr_09x_01)));
      state_10( 6) <= S_BOX_10_06(to_integer(unsigned(addr_09x_01)));
      state_10( 7) <= S_BOX_10_07(to_integer(unsigned(addr_09x_01)));
      state_10( 8) <= S_BOX_10_08(to_integer(unsigned(addr_09x_02)));
      state_10( 9) <= S_BOX_10_09(to_integer(unsigned(addr_09x_02)));
      state_10(10) <= S_BOX_10_10(to_integer(unsigned(addr_09x_02)));
      state_10(11) <= S_BOX_10_11(to_integer(unsigned(addr_09x_02)));
      state_10(12) <= S_BOX_10_12(to_integer(unsigned(addr_09x_03)));
      state_10(13) <= S_BOX_10_13(to_integer(unsigned(addr_09x_03)));
      state_10(14) <= S_BOX_10_14(to_integer(unsigned(addr_09x_03)));
      state_10(15) <= S_BOX_10_15(to_integer(unsigned(addr_09x_03)));
      state_10(16) <= S_BOX_10_16(to_integer(unsigned(addr_09x_04)));
      state_10(17) <= S_BOX_10_17(to_integer(unsigned(addr_09x_04)));
      state_10(18) <= S_BOX_10_18(to_integer(unsigned(addr_09x_04)));
      state_10(19) <= S_BOX_10_19(to_integer(unsigned(addr_09x_04)));
      state_10(20) <= S_BOX_10_20(to_integer(unsigned(addr_09x_05)));
      state_10(21) <= S_BOX_10_21(to_integer(unsigned(addr_09x_05)));
      state_10(22) <= S_BOX_10_22(to_integer(unsigned(addr_09x_05)));
      state_10(23) <= S_BOX_10_23(to_integer(unsigned(addr_09x_05)));
      state_10(24) <= S_BOX_10_24(to_integer(unsigned(addr_09x_06)));
      state_10(25) <= S_BOX_10_25(to_integer(unsigned(addr_09x_06)));
      state_10(26) <= S_BOX_10_26(to_integer(unsigned(addr_09x_06)));
      state_10(27) <= S_BOX_10_27(to_integer(unsigned(addr_09x_06)));
      state_10(28) <= S_BOX_10_28(to_integer(unsigned(addr_09x_07)));
      state_10(29) <= S_BOX_10_29(to_integer(unsigned(addr_09x_07)));
      state_10(30) <= S_BOX_10_30(to_integer(unsigned(addr_09x_07)));
      state_10(31) <= S_BOX_10_31(to_integer(unsigned(addr_09x_07)));
      state_10(32) <= S_BOX_10_32(to_integer(unsigned(addr_09x_08)));
      state_10(33) <= S_BOX_10_33(to_integer(unsigned(addr_09x_08)));
      state_10(34) <= S_BOX_10_34(to_integer(unsigned(addr_09x_08)));
      state_10(35) <= S_BOX_10_35(to_integer(unsigned(addr_09x_08)));
      state_10(36) <= S_BOX_10_36(to_integer(unsigned(addr_09x_09)));
      state_10(37) <= S_BOX_10_37(to_integer(unsigned(addr_09x_09)));
      state_10(38) <= S_BOX_10_38(to_integer(unsigned(addr_09x_09)));
      state_10(39) <= S_BOX_10_39(to_integer(unsigned(addr_09x_09)));
      state_10(40) <= S_BOX_10_40(to_integer(unsigned(addr_09x_10)));
      state_10(41) <= S_BOX_10_41(to_integer(unsigned(addr_09x_10)));
      state_10(42) <= S_BOX_10_42(to_integer(unsigned(addr_09x_10)));
      state_10(43) <= S_BOX_10_43(to_integer(unsigned(addr_09x_10)));
      state_10(44) <= S_BOX_10_44(to_integer(unsigned(addr_09x_11)));
      state_10(45) <= S_BOX_10_45(to_integer(unsigned(addr_09x_11)));
      state_10(46) <= S_BOX_10_46(to_integer(unsigned(addr_09x_11)));
      state_10(47) <= S_BOX_10_47(to_integer(unsigned(addr_09x_11)));
    end if;
  end process;
end heavy;

--
-- Warped linear feedback shift register pseudo-random number generator (period=2^48-1)
--
architecture light of pseudo_random_generator is
  constant ZERO       : std_logic_vector(47 downto 0) := (others => '0'); -- the zero constant
  signal   state      : std_logic_vector(47 downto 0) := SEED;            -- the current pseudo-random generator state
  signal   next_state : std_logic_vector(47 downto 0);                    -- the next pseudo-random generator state
  signal   kick       : std_logic;                                        -- set to one if the state is zero
begin
  --
  -- Output
  --
  rnd <= state(N_BITS-1 downto 0);
  --
  -- State update
  --
  process(enable,clock) is
  begin
    if enable = '1' and rising_edge(clock) then
      if state = ZERO then -- this can only happen if SEED = ZERO or if there is a hardware error
        kick <= '1';
      else
        kick <= '0';
      end if;
      state <= next_state;
    end if;
  end process;
  --
  -- Next state computation (data generated by c_code/pseudo_random_generator.c with n=48 and seed=1)
  --
  next_state( 0) <= state(17) xor state(27) xor state(30) xor state(33); -- state( 0) used  5 times
  next_state( 1) <= state(21) xor state(28) xor state(29) xor kick;      -- state( 1) used  2 times
  next_state( 2) <= state( 8) xor state(22) xor state(33) xor state(35); -- state( 2) used  2 times
  next_state( 3) <= state( 9) xor state(14) xor state(21) xor state(47); -- state( 3) used  5 times
  next_state( 4) <= state( 3) xor state(24) xor state(32) xor state(44); -- state( 4) used  2 times
  next_state( 5) <= state(10) xor state(15) xor state(27) xor state(44); -- state( 5) used  4 times
  next_state( 6) <= state( 7) xor state(10) xor state(16) xor state(46); -- state( 6) used  4 times
  next_state( 7) <= state(25) xor state(27) xor state(28) xor state(31); -- state( 7) used  5 times
  next_state( 8) <= state( 2) xor state(17) xor state(25) xor state(31); -- state( 8) used  4 times
  next_state( 9) <= state(12) xor state(24) xor state(35);               -- state( 9) used  4 times
  next_state(10) <= state(10) xor state(14) xor state(16) xor state(22); -- state(10) used  5 times
  next_state(11) <= state( 5) xor state(18) xor state(35) xor state(47); -- state(11) used  2 times
  next_state(12) <= state(19) xor state(28) xor state(31) xor state(45); -- state(12) used  3 times
  next_state(13) <= state(23) xor state(37) xor state(40) xor state(43); -- state(13) used  5 times
  next_state(14) <= state(21) xor state(30) xor state(32) xor state(42); -- state(14) used  2 times
  next_state(15) <= state( 3) xor state( 5) xor state(39) xor state(40); -- state(15) used  2 times
  next_state(16) <= state( 0) xor state(29) xor state(37) xor state(45); -- state(16) used  5 times
  next_state(17) <= state( 4) xor state(26) xor state(38) xor state(47); -- state(17) used  5 times
  next_state(18) <= state( 8) xor state(13) xor state(40) xor state(42); -- state(18) used  5 times
  next_state(19) <= state(20) xor state(32) xor state(35) xor state(38); -- state(19) used  3 times
  next_state(20) <= state(11) xor state(33) xor state(39) xor state(45); -- state(20) used  5 times
  next_state(21) <= state(16) xor state(18) xor state(24) xor state(35); -- state(21) used  5 times
  next_state(22) <= state( 0) xor state(34) xor state(38) xor state(42); -- state(22) used  2 times
  next_state(23) <= state(20) xor state(21) xor state(40) xor state(46); -- state(23) used  2 times
  next_state(24) <= state(18) xor state(28) xor state(31) xor state(34); -- state(24) used  3 times
  next_state(25) <= state(11) xor state(18) xor state(20) xor state(44); -- state(25) used  5 times
  next_state(26) <= state(19) xor state(29) xor state(33) xor state(45); -- state(26) used  3 times
  next_state(27) <= state( 3) xor state(16) xor state(26) xor state(34); -- state(27) used  4 times
  next_state(28) <= state( 8) xor state(15) xor state(17) xor state(20); -- state(28) used  5 times
  next_state(29) <= state( 6) xor state( 8) xor state(25) xor state(36); -- state(29) used  5 times
  next_state(30) <= state(13) xor state(17) xor state(25) xor state(34); -- state(30) used  5 times
  next_state(31) <= state(10) xor state(33) xor state(34) xor state(44); -- state(31) used  5 times
  next_state(32) <= state( 9) xor state(12) xor state(17) xor state(21); -- state(32) used  4 times
  next_state(33) <= state( 5) xor state( 6) xor state(30) xor state(41); -- state(33) used  5 times
  next_state(34) <= state( 0) xor state(13) xor state(25) xor state(38); -- state(34) used  5 times
  next_state(35) <= state( 3) xor state(16) xor state(18) xor state(36); -- state(35) used  5 times
  next_state(36) <= state( 6) xor state(28) xor state(37) xor state(41); -- state(36) used  4 times
  next_state(37) <= state( 0) xor state( 1) xor state(13) xor state(45); -- state(37) used  5 times
  next_state(38) <= state(29) xor state(31) xor state(36) xor state(46); -- state(38) used  4 times
  next_state(39) <= state( 2) xor state( 6) xor state( 7) xor state(37); -- state(39) used  3 times
  next_state(40) <= state(23) xor state(26) xor state(37) xor state(46); -- state(40) used  5 times
  next_state(41) <= state(13) xor state(19) xor state(20) xor state(43); -- state(41) used  2 times
  next_state(42) <= state( 5) xor state( 7) xor state(12) xor state(29); -- state(42) used  5 times
  next_state(43) <= state( 9) xor state(30) xor state(40) xor state(42); -- state(43) used  2 times
  next_state(44) <= state( 4) xor state( 7) xor state(30) xor state(44); -- state(44) used  5 times
  next_state(45) <= state( 1) xor state( 3) xor state( 7) xor state(46); -- state(45) used  5 times
  next_state(46) <= state(27) xor state(32) xor state(39) xor state(42); -- state(46) used  5 times
  next_state(47) <= state( 0) xor state( 9) xor state(10) xor state(36); -- state(47) used  3 times
end light;
